// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : PoseidonTopLevel


`define ReceiverState_binary_sequential_type [2:0]
`define ReceiverState_binary_sequential_IDLE 3'b000
`define ReceiverState_binary_sequential_ELEMENT0 3'b001
`define ReceiverState_binary_sequential_ELEMENT1 3'b010
`define ReceiverState_binary_sequential_BLOCK_1 3'b011
`define ReceiverState_binary_sequential_BLOCK_IDLE 3'b100
`define ReceiverState_binary_sequential_DONE 3'b101

`define threadAccumulator_fsm_enumDefinition_binary_sequential_type [1:0]
`define threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_BOOT 2'b00
`define threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE 2'b01
`define threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING 2'b10
`define threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE 2'b11


module PoseidonTopLevel (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_last,
  input      [254:0]  io_input_payload,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_last,
  output     [254:0]  io_output_payload,
  input               reset,
  input               clk
);
  wire                receiver_io_outputs_0_ready;
  wire                receiver_io_outputs_1_ready;
  wire                receiver_io_outputs_2_ready;
  wire                receiver_io_input_ready;
  wire                receiver_io_outputs_0_valid;
  wire       [6:0]    receiver_io_outputs_0_payload_round_index;
  wire       [3:0]    receiver_io_outputs_0_payload_state_index;
  wire       [3:0]    receiver_io_outputs_0_payload_state_size;
  wire       [6:0]    receiver_io_outputs_0_payload_state_id;
  wire       [254:0]  receiver_io_outputs_0_payload_state_element;
  wire                receiver_io_outputs_1_valid;
  wire       [6:0]    receiver_io_outputs_1_payload_round_index;
  wire       [3:0]    receiver_io_outputs_1_payload_state_index;
  wire       [3:0]    receiver_io_outputs_1_payload_state_size;
  wire       [6:0]    receiver_io_outputs_1_payload_state_id;
  wire       [254:0]  receiver_io_outputs_1_payload_state_element;
  wire                receiver_io_outputs_2_valid;
  wire       [6:0]    receiver_io_outputs_2_payload_round_index;
  wire       [3:0]    receiver_io_outputs_2_payload_state_index;
  wire       [3:0]    receiver_io_outputs_2_payload_state_size;
  wire       [6:0]    receiver_io_outputs_2_payload_state_id;
  wire       [254:0]  receiver_io_outputs_2_payload_state_element;
  wire                streamArbiter_12_io_inputs_0_ready;
  wire                streamArbiter_12_io_inputs_1_ready;
  wire                streamArbiter_12_io_output_valid;
  wire       [6:0]    streamArbiter_12_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_12_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_12_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_12_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_12_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_12_io_chosen;
  wire       [1:0]    streamArbiter_12_io_chosenOH;
  wire                streamArbiter_13_io_inputs_0_ready;
  wire                streamArbiter_13_io_inputs_1_ready;
  wire                streamArbiter_13_io_output_valid;
  wire       [6:0]    streamArbiter_13_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_13_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_13_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_13_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_13_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_13_io_chosen;
  wire       [1:0]    streamArbiter_13_io_chosenOH;
  wire                streamArbiter_14_io_inputs_0_ready;
  wire                streamArbiter_14_io_inputs_1_ready;
  wire                streamArbiter_14_io_output_valid;
  wire       [6:0]    streamArbiter_14_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_14_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_14_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_14_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_14_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_14_io_chosen;
  wire       [1:0]    streamArbiter_14_io_chosenOH;
  wire                DataProcess_matrixAdder_io_inputs_0_ready;
  wire                DataProcess_matrixAdder_io_inputs_1_ready;
  wire                DataProcess_matrixAdder_io_inputs_2_ready;
  wire                DataProcess_matrixAdder_io_output_valid;
  wire       [6:0]    DataProcess_matrixAdder_io_output_payload_round_index;
  wire       [3:0]    DataProcess_matrixAdder_io_output_payload_state_size;
  wire       [6:0]    DataProcess_matrixAdder_io_output_payload_state_id;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_0;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_1;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_2;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_3;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_4;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_5;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_6;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_7;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_8;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_9;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_10;
  wire       [254:0]  DataProcess_matrixAdder_io_output_payload_state_elements_11;
  wire                poseidonThread_3_io_input_ready;
  wire                poseidonThread_3_io_output_valid;
  wire       [6:0]    poseidonThread_3_io_output_payload_round_index;
  wire       [3:0]    poseidonThread_3_io_output_payload_state_size;
  wire       [6:0]    poseidonThread_3_io_output_payload_state_id;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_0;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_1;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_2;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_3;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_4;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_5;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_6;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_7;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_8;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_9;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_10;
  wire       [254:0]  poseidonThread_3_io_output_payload_state_elements_11;
  wire                poseidonThread_4_io_input_ready;
  wire                poseidonThread_4_io_output_valid;
  wire       [6:0]    poseidonThread_4_io_output_payload_round_index;
  wire       [3:0]    poseidonThread_4_io_output_payload_state_size;
  wire       [6:0]    poseidonThread_4_io_output_payload_state_id;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_0;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_1;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_2;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_3;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_4;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_5;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_6;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_7;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_8;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_9;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_10;
  wire       [254:0]  poseidonThread_4_io_output_payload_state_elements_11;
  wire                poseidonThread_5_io_input_ready;
  wire                poseidonThread_5_io_output_valid;
  wire       [6:0]    poseidonThread_5_io_output_payload_round_index;
  wire       [3:0]    poseidonThread_5_io_output_payload_state_size;
  wire       [6:0]    poseidonThread_5_io_output_payload_state_id;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_0;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_1;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_2;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_3;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_4;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_5;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_6;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_7;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_8;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_9;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_10;
  wire       [254:0]  poseidonThread_5_io_output_payload_state_elements_11;
  wire                loopbackBuffer_io_input_ready;
  wire                loopbackBuffer_io_outputs_0_valid;
  wire       [6:0]    loopbackBuffer_io_outputs_0_payload_round_index;
  wire       [3:0]    loopbackBuffer_io_outputs_0_payload_state_index;
  wire       [3:0]    loopbackBuffer_io_outputs_0_payload_state_size;
  wire       [6:0]    loopbackBuffer_io_outputs_0_payload_state_id;
  wire       [254:0]  loopbackBuffer_io_outputs_0_payload_state_element;
  wire                loopbackBuffer_io_outputs_1_valid;
  wire       [6:0]    loopbackBuffer_io_outputs_1_payload_round_index;
  wire       [3:0]    loopbackBuffer_io_outputs_1_payload_state_index;
  wire       [3:0]    loopbackBuffer_io_outputs_1_payload_state_size;
  wire       [6:0]    loopbackBuffer_io_outputs_1_payload_state_id;
  wire       [254:0]  loopbackBuffer_io_outputs_1_payload_state_element;
  wire                loopbackBuffer_io_outputs_2_valid;
  wire       [6:0]    loopbackBuffer_io_outputs_2_payload_round_index;
  wire       [3:0]    loopbackBuffer_io_outputs_2_payload_state_index;
  wire       [3:0]    loopbackBuffer_io_outputs_2_payload_state_size;
  wire       [6:0]    loopbackBuffer_io_outputs_2_payload_state_id;
  wire       [254:0]  loopbackBuffer_io_outputs_2_payload_state_element;
  wire       [3:0]    loopbackBuffer_io_residue;
  wire                transmitter_io_input_ready;
  wire                transmitter_io_output_valid;
  wire                transmitter_io_output_last;
  wire       [254:0]  transmitter_io_output_payload;
  wire       [3:0]    _zz__zz_DataMux_inputs1_temp_0_ready;
  wire       [3:0]    _zz__zz_DataMux_inputs1_temp_1_ready;
  wire       [3:0]    _zz__zz_DataMux_inputs1_temp_2_ready;
  wire                DataMux_inputs0_0_valid;
  wire                DataMux_inputs0_0_ready;
  wire       [6:0]    DataMux_inputs0_0_payload_round_index;
  wire       [3:0]    DataMux_inputs0_0_payload_state_index;
  wire       [3:0]    DataMux_inputs0_0_payload_state_size;
  wire       [6:0]    DataMux_inputs0_0_payload_state_id;
  wire       [254:0]  DataMux_inputs0_0_payload_state_element;
  wire                DataMux_inputs0_1_valid;
  wire                DataMux_inputs0_1_ready;
  wire       [6:0]    DataMux_inputs0_1_payload_round_index;
  wire       [3:0]    DataMux_inputs0_1_payload_state_index;
  wire       [3:0]    DataMux_inputs0_1_payload_state_size;
  wire       [6:0]    DataMux_inputs0_1_payload_state_id;
  wire       [254:0]  DataMux_inputs0_1_payload_state_element;
  wire                DataMux_inputs0_2_valid;
  wire                DataMux_inputs0_2_ready;
  wire       [6:0]    DataMux_inputs0_2_payload_round_index;
  wire       [3:0]    DataMux_inputs0_2_payload_state_index;
  wire       [3:0]    DataMux_inputs0_2_payload_state_size;
  wire       [6:0]    DataMux_inputs0_2_payload_state_id;
  wire       [254:0]  DataMux_inputs0_2_payload_state_element;
  wire                DataMux_inputs1_temp_0_valid;
  wire                DataMux_inputs1_temp_0_ready;
  wire       [6:0]    DataMux_inputs1_temp_0_payload_round_index;
  wire       [3:0]    DataMux_inputs1_temp_0_payload_state_index;
  wire       [3:0]    DataMux_inputs1_temp_0_payload_state_size;
  wire       [6:0]    DataMux_inputs1_temp_0_payload_state_id;
  wire       [254:0]  DataMux_inputs1_temp_0_payload_state_element;
  wire                DataMux_inputs1_temp_1_valid;
  wire                DataMux_inputs1_temp_1_ready;
  wire       [6:0]    DataMux_inputs1_temp_1_payload_round_index;
  wire       [3:0]    DataMux_inputs1_temp_1_payload_state_index;
  wire       [3:0]    DataMux_inputs1_temp_1_payload_state_size;
  wire       [6:0]    DataMux_inputs1_temp_1_payload_state_id;
  wire       [254:0]  DataMux_inputs1_temp_1_payload_state_element;
  wire                DataMux_inputs1_temp_2_valid;
  wire                DataMux_inputs1_temp_2_ready;
  wire       [6:0]    DataMux_inputs1_temp_2_payload_round_index;
  wire       [3:0]    DataMux_inputs1_temp_2_payload_state_index;
  wire       [3:0]    DataMux_inputs1_temp_2_payload_state_size;
  wire       [6:0]    DataMux_inputs1_temp_2_payload_state_id;
  wire       [254:0]  DataMux_inputs1_temp_2_payload_state_element;
  wire                receiver_io_outputs_0_s2mPipe_valid;
  reg                 receiver_io_outputs_0_s2mPipe_ready;
  wire       [6:0]    receiver_io_outputs_0_s2mPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_0_s2mPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_0_s2mPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_0_s2mPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_0_s2mPipe_payload_state_element;
  reg                 receiver_io_outputs_0_rValid;
  reg        [6:0]    receiver_io_outputs_0_rData_round_index;
  reg        [3:0]    receiver_io_outputs_0_rData_state_index;
  reg        [3:0]    receiver_io_outputs_0_rData_state_size;
  reg        [6:0]    receiver_io_outputs_0_rData_state_id;
  reg        [254:0]  receiver_io_outputs_0_rData_state_element;
  wire                receiver_io_outputs_0_s2mPipe_m2sPipe_valid;
  wire                receiver_io_outputs_0_s2mPipe_m2sPipe_ready;
  wire       [6:0]    receiver_io_outputs_0_s2mPipe_m2sPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_element;
  reg                 receiver_io_outputs_0_s2mPipe_rValid;
  reg        [6:0]    receiver_io_outputs_0_s2mPipe_rData_round_index;
  reg        [3:0]    receiver_io_outputs_0_s2mPipe_rData_state_index;
  reg        [3:0]    receiver_io_outputs_0_s2mPipe_rData_state_size;
  reg        [6:0]    receiver_io_outputs_0_s2mPipe_rData_state_id;
  reg        [254:0]  receiver_io_outputs_0_s2mPipe_rData_state_element;
  wire                when_Stream_l342;
  wire                receiver_io_outputs_1_s2mPipe_valid;
  reg                 receiver_io_outputs_1_s2mPipe_ready;
  wire       [6:0]    receiver_io_outputs_1_s2mPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_1_s2mPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_1_s2mPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_1_s2mPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_1_s2mPipe_payload_state_element;
  reg                 receiver_io_outputs_1_rValid;
  reg        [6:0]    receiver_io_outputs_1_rData_round_index;
  reg        [3:0]    receiver_io_outputs_1_rData_state_index;
  reg        [3:0]    receiver_io_outputs_1_rData_state_size;
  reg        [6:0]    receiver_io_outputs_1_rData_state_id;
  reg        [254:0]  receiver_io_outputs_1_rData_state_element;
  wire                receiver_io_outputs_1_s2mPipe_m2sPipe_valid;
  wire                receiver_io_outputs_1_s2mPipe_m2sPipe_ready;
  wire       [6:0]    receiver_io_outputs_1_s2mPipe_m2sPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_element;
  reg                 receiver_io_outputs_1_s2mPipe_rValid;
  reg        [6:0]    receiver_io_outputs_1_s2mPipe_rData_round_index;
  reg        [3:0]    receiver_io_outputs_1_s2mPipe_rData_state_index;
  reg        [3:0]    receiver_io_outputs_1_s2mPipe_rData_state_size;
  reg        [6:0]    receiver_io_outputs_1_s2mPipe_rData_state_id;
  reg        [254:0]  receiver_io_outputs_1_s2mPipe_rData_state_element;
  wire                when_Stream_l342_1;
  wire                receiver_io_outputs_2_s2mPipe_valid;
  reg                 receiver_io_outputs_2_s2mPipe_ready;
  wire       [6:0]    receiver_io_outputs_2_s2mPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_2_s2mPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_2_s2mPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_2_s2mPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_2_s2mPipe_payload_state_element;
  reg                 receiver_io_outputs_2_rValid;
  reg        [6:0]    receiver_io_outputs_2_rData_round_index;
  reg        [3:0]    receiver_io_outputs_2_rData_state_index;
  reg        [3:0]    receiver_io_outputs_2_rData_state_size;
  reg        [6:0]    receiver_io_outputs_2_rData_state_id;
  reg        [254:0]  receiver_io_outputs_2_rData_state_element;
  wire                receiver_io_outputs_2_s2mPipe_m2sPipe_valid;
  wire                receiver_io_outputs_2_s2mPipe_m2sPipe_ready;
  wire       [6:0]    receiver_io_outputs_2_s2mPipe_m2sPipe_payload_round_index;
  wire       [3:0]    receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_index;
  wire       [3:0]    receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_size;
  wire       [6:0]    receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_id;
  wire       [254:0]  receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_element;
  reg                 receiver_io_outputs_2_s2mPipe_rValid;
  reg        [6:0]    receiver_io_outputs_2_s2mPipe_rData_round_index;
  reg        [3:0]    receiver_io_outputs_2_s2mPipe_rData_state_index;
  reg        [3:0]    receiver_io_outputs_2_s2mPipe_rData_state_size;
  reg        [6:0]    receiver_io_outputs_2_s2mPipe_rData_state_id;
  reg        [254:0]  receiver_io_outputs_2_s2mPipe_rData_state_element;
  wire                when_Stream_l342_2;
  wire       [3:0]    DataMux_residue;
  wire                _zz_DataMux_inputs1_temp_0_ready;
  wire                DataMux_inputs1_0_valid;
  wire                DataMux_inputs1_0_ready;
  wire       [6:0]    DataMux_inputs1_0_payload_round_index;
  wire       [3:0]    DataMux_inputs1_0_payload_state_index;
  wire       [3:0]    DataMux_inputs1_0_payload_state_size;
  wire       [6:0]    DataMux_inputs1_0_payload_state_id;
  wire       [254:0]  DataMux_inputs1_0_payload_state_element;
  wire                _zz_DataMux_inputs1_temp_1_ready;
  wire                DataMux_inputs1_1_valid;
  wire                DataMux_inputs1_1_ready;
  wire       [6:0]    DataMux_inputs1_1_payload_round_index;
  wire       [3:0]    DataMux_inputs1_1_payload_state_index;
  wire       [3:0]    DataMux_inputs1_1_payload_state_size;
  wire       [6:0]    DataMux_inputs1_1_payload_state_id;
  wire       [254:0]  DataMux_inputs1_1_payload_state_element;
  wire                _zz_DataMux_inputs1_temp_2_ready;
  wire                DataMux_inputs1_2_valid;
  wire                DataMux_inputs1_2_ready;
  wire       [6:0]    DataMux_inputs1_2_payload_round_index;
  wire       [3:0]    DataMux_inputs1_2_payload_state_index;
  wire       [3:0]    DataMux_inputs1_2_payload_state_size;
  wire       [6:0]    DataMux_inputs1_2_payload_state_id;
  wire       [254:0]  DataMux_inputs1_2_payload_state_element;
  wire                DataMux_outputs_0_valid;
  wire                DataMux_outputs_0_ready;
  wire       [6:0]    DataMux_outputs_0_payload_round_index;
  wire       [3:0]    DataMux_outputs_0_payload_state_index;
  wire       [3:0]    DataMux_outputs_0_payload_state_size;
  wire       [6:0]    DataMux_outputs_0_payload_state_id;
  wire       [254:0]  DataMux_outputs_0_payload_state_element;
  wire                DataMux_outputs_1_valid;
  wire                DataMux_outputs_1_ready;
  wire       [6:0]    DataMux_outputs_1_payload_round_index;
  wire       [3:0]    DataMux_outputs_1_payload_state_index;
  wire       [3:0]    DataMux_outputs_1_payload_state_size;
  wire       [6:0]    DataMux_outputs_1_payload_state_id;
  wire       [254:0]  DataMux_outputs_1_payload_state_element;
  wire                DataMux_outputs_2_valid;
  wire                DataMux_outputs_2_ready;
  wire       [6:0]    DataMux_outputs_2_payload_round_index;
  wire       [3:0]    DataMux_outputs_2_payload_state_index;
  wire       [3:0]    DataMux_outputs_2_payload_state_size;
  wire       [6:0]    DataMux_outputs_2_payload_state_id;
  wire       [254:0]  DataMux_outputs_2_payload_state_element;
  wire                DataProcess_output_valid;
  wire                DataProcess_output_ready;
  wire       [6:0]    DataProcess_output_payload_round_index;
  wire       [3:0]    DataProcess_output_payload_state_size;
  wire       [6:0]    DataProcess_output_payload_state_id;
  wire       [254:0]  DataProcess_output_payload_state_elements_0;
  wire       [254:0]  DataProcess_output_payload_state_elements_1;
  wire       [254:0]  DataProcess_output_payload_state_elements_2;
  wire       [254:0]  DataProcess_output_payload_state_elements_3;
  wire       [254:0]  DataProcess_output_payload_state_elements_4;
  wire       [254:0]  DataProcess_output_payload_state_elements_5;
  wire       [254:0]  DataProcess_output_payload_state_elements_6;
  wire       [254:0]  DataProcess_output_payload_state_elements_7;
  wire       [254:0]  DataProcess_output_payload_state_elements_8;
  wire       [254:0]  DataProcess_output_payload_state_elements_9;
  wire       [254:0]  DataProcess_output_payload_state_elements_10;
  wire       [254:0]  DataProcess_output_payload_state_elements_11;
  wire                DataDeMux_output0_valid;
  wire                DataDeMux_output0_ready;
  wire       [6:0]    DataDeMux_output0_payload_state_id;
  wire       [254:0]  DataDeMux_output0_payload_state_element;
  wire                DataDeMux_output1_valid;
  wire                DataDeMux_output1_ready;
  reg        [6:0]    DataDeMux_output1_payload_round_index;
  wire       [3:0]    DataDeMux_output1_payload_state_size;
  wire       [6:0]    DataDeMux_output1_payload_state_id;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_0;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_1;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_2;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_3;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_4;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_5;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_6;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_7;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_8;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_9;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_10;
  wire       [254:0]  DataDeMux_output1_payload_state_elements_11;
  reg        [1:0]    DataDeMux_select;

  assign _zz__zz_DataMux_inputs1_temp_0_ready = (DataMux_inputs1_temp_0_payload_state_size - DataMux_inputs1_temp_0_payload_state_index);
  assign _zz__zz_DataMux_inputs1_temp_1_ready = (DataMux_inputs1_temp_0_payload_state_size - DataMux_inputs1_temp_0_payload_state_index);
  assign _zz__zz_DataMux_inputs1_temp_2_ready = (DataMux_inputs1_temp_0_payload_state_size - DataMux_inputs1_temp_0_payload_state_index);
  AXI4StreamReceiver receiver (
    .io_input_valid                        (io_input_valid                               ), //i
    .io_input_ready                        (receiver_io_input_ready                      ), //o
    .io_input_last                         (io_input_last                                ), //i
    .io_input_payload                      (io_input_payload                             ), //i
    .io_outputs_0_valid                    (receiver_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (receiver_io_outputs_0_ready                  ), //i
    .io_outputs_0_payload_round_index      (receiver_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (receiver_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (receiver_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (receiver_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (receiver_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (receiver_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (receiver_io_outputs_1_ready                  ), //i
    .io_outputs_1_payload_round_index      (receiver_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (receiver_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (receiver_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (receiver_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (receiver_io_outputs_1_payload_state_element  ), //o
    .io_outputs_2_valid                    (receiver_io_outputs_2_valid                  ), //o
    .io_outputs_2_ready                    (receiver_io_outputs_2_ready                  ), //i
    .io_outputs_2_payload_round_index      (receiver_io_outputs_2_payload_round_index    ), //o
    .io_outputs_2_payload_state_index      (receiver_io_outputs_2_payload_state_index    ), //o
    .io_outputs_2_payload_state_size       (receiver_io_outputs_2_payload_state_size     ), //o
    .io_outputs_2_payload_state_id         (receiver_io_outputs_2_payload_state_id       ), //o
    .io_outputs_2_payload_state_element    (receiver_io_outputs_2_payload_state_element  ), //o
    .clk                                   (clk                                          ), //i
    .reset                                 (reset                                        )  //i
  );
  StreamArbiter streamArbiter_12 (
    .io_inputs_0_valid                    (DataMux_inputs0_0_valid                           ), //i
    .io_inputs_0_ready                    (streamArbiter_12_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (DataMux_inputs0_0_payload_round_index             ), //i
    .io_inputs_0_payload_state_index      (DataMux_inputs0_0_payload_state_index             ), //i
    .io_inputs_0_payload_state_size       (DataMux_inputs0_0_payload_state_size              ), //i
    .io_inputs_0_payload_state_id         (DataMux_inputs0_0_payload_state_id                ), //i
    .io_inputs_0_payload_state_element    (DataMux_inputs0_0_payload_state_element           ), //i
    .io_inputs_1_valid                    (DataMux_inputs1_0_valid                           ), //i
    .io_inputs_1_ready                    (streamArbiter_12_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (DataMux_inputs1_0_payload_round_index             ), //i
    .io_inputs_1_payload_state_index      (DataMux_inputs1_0_payload_state_index             ), //i
    .io_inputs_1_payload_state_size       (DataMux_inputs1_0_payload_state_size              ), //i
    .io_inputs_1_payload_state_id         (DataMux_inputs1_0_payload_state_id                ), //i
    .io_inputs_1_payload_state_element    (DataMux_inputs1_0_payload_state_element           ), //i
    .io_output_valid                      (streamArbiter_12_io_output_valid                  ), //o
    .io_output_ready                      (DataMux_outputs_0_ready                           ), //i
    .io_output_payload_round_index        (streamArbiter_12_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_12_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_12_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_12_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_12_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_12_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_12_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_13 (
    .io_inputs_0_valid                    (DataMux_inputs0_1_valid                           ), //i
    .io_inputs_0_ready                    (streamArbiter_13_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (DataMux_inputs0_1_payload_round_index             ), //i
    .io_inputs_0_payload_state_index      (DataMux_inputs0_1_payload_state_index             ), //i
    .io_inputs_0_payload_state_size       (DataMux_inputs0_1_payload_state_size              ), //i
    .io_inputs_0_payload_state_id         (DataMux_inputs0_1_payload_state_id                ), //i
    .io_inputs_0_payload_state_element    (DataMux_inputs0_1_payload_state_element           ), //i
    .io_inputs_1_valid                    (DataMux_inputs1_1_valid                           ), //i
    .io_inputs_1_ready                    (streamArbiter_13_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (DataMux_inputs1_1_payload_round_index             ), //i
    .io_inputs_1_payload_state_index      (DataMux_inputs1_1_payload_state_index             ), //i
    .io_inputs_1_payload_state_size       (DataMux_inputs1_1_payload_state_size              ), //i
    .io_inputs_1_payload_state_id         (DataMux_inputs1_1_payload_state_id                ), //i
    .io_inputs_1_payload_state_element    (DataMux_inputs1_1_payload_state_element           ), //i
    .io_output_valid                      (streamArbiter_13_io_output_valid                  ), //o
    .io_output_ready                      (DataMux_outputs_1_ready                           ), //i
    .io_output_payload_round_index        (streamArbiter_13_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_13_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_13_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_13_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_13_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_13_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_13_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_14 (
    .io_inputs_0_valid                    (DataMux_inputs0_2_valid                           ), //i
    .io_inputs_0_ready                    (streamArbiter_14_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (DataMux_inputs0_2_payload_round_index             ), //i
    .io_inputs_0_payload_state_index      (DataMux_inputs0_2_payload_state_index             ), //i
    .io_inputs_0_payload_state_size       (DataMux_inputs0_2_payload_state_size              ), //i
    .io_inputs_0_payload_state_id         (DataMux_inputs0_2_payload_state_id                ), //i
    .io_inputs_0_payload_state_element    (DataMux_inputs0_2_payload_state_element           ), //i
    .io_inputs_1_valid                    (DataMux_inputs1_2_valid                           ), //i
    .io_inputs_1_ready                    (streamArbiter_14_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (DataMux_inputs1_2_payload_round_index             ), //i
    .io_inputs_1_payload_state_index      (DataMux_inputs1_2_payload_state_index             ), //i
    .io_inputs_1_payload_state_size       (DataMux_inputs1_2_payload_state_size              ), //i
    .io_inputs_1_payload_state_id         (DataMux_inputs1_2_payload_state_id                ), //i
    .io_inputs_1_payload_state_element    (DataMux_inputs1_2_payload_state_element           ), //i
    .io_output_valid                      (streamArbiter_14_io_output_valid                  ), //o
    .io_output_ready                      (DataMux_outputs_2_ready                           ), //i
    .io_output_payload_round_index        (streamArbiter_14_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_14_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_14_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_14_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_14_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_14_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_14_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  MDSMatrixAdders DataProcess_matrixAdder (
    .io_inputs_0_valid                        (poseidonThread_3_io_output_valid                             ), //i
    .io_inputs_0_ready                        (DataProcess_matrixAdder_io_inputs_0_ready                    ), //o
    .io_inputs_0_payload_round_index          (poseidonThread_3_io_output_payload_round_index               ), //i
    .io_inputs_0_payload_state_size           (poseidonThread_3_io_output_payload_state_size                ), //i
    .io_inputs_0_payload_state_id             (poseidonThread_3_io_output_payload_state_id                  ), //i
    .io_inputs_0_payload_state_elements_0     (poseidonThread_3_io_output_payload_state_elements_0          ), //i
    .io_inputs_0_payload_state_elements_1     (poseidonThread_3_io_output_payload_state_elements_1          ), //i
    .io_inputs_0_payload_state_elements_2     (poseidonThread_3_io_output_payload_state_elements_2          ), //i
    .io_inputs_0_payload_state_elements_3     (poseidonThread_3_io_output_payload_state_elements_3          ), //i
    .io_inputs_0_payload_state_elements_4     (poseidonThread_3_io_output_payload_state_elements_4          ), //i
    .io_inputs_0_payload_state_elements_5     (poseidonThread_3_io_output_payload_state_elements_5          ), //i
    .io_inputs_0_payload_state_elements_6     (poseidonThread_3_io_output_payload_state_elements_6          ), //i
    .io_inputs_0_payload_state_elements_7     (poseidonThread_3_io_output_payload_state_elements_7          ), //i
    .io_inputs_0_payload_state_elements_8     (poseidonThread_3_io_output_payload_state_elements_8          ), //i
    .io_inputs_0_payload_state_elements_9     (poseidonThread_3_io_output_payload_state_elements_9          ), //i
    .io_inputs_0_payload_state_elements_10    (poseidonThread_3_io_output_payload_state_elements_10         ), //i
    .io_inputs_0_payload_state_elements_11    (poseidonThread_3_io_output_payload_state_elements_11         ), //i
    .io_inputs_1_valid                        (poseidonThread_4_io_output_valid                             ), //i
    .io_inputs_1_ready                        (DataProcess_matrixAdder_io_inputs_1_ready                    ), //o
    .io_inputs_1_payload_round_index          (poseidonThread_4_io_output_payload_round_index               ), //i
    .io_inputs_1_payload_state_size           (poseidonThread_4_io_output_payload_state_size                ), //i
    .io_inputs_1_payload_state_id             (poseidonThread_4_io_output_payload_state_id                  ), //i
    .io_inputs_1_payload_state_elements_0     (poseidonThread_4_io_output_payload_state_elements_0          ), //i
    .io_inputs_1_payload_state_elements_1     (poseidonThread_4_io_output_payload_state_elements_1          ), //i
    .io_inputs_1_payload_state_elements_2     (poseidonThread_4_io_output_payload_state_elements_2          ), //i
    .io_inputs_1_payload_state_elements_3     (poseidonThread_4_io_output_payload_state_elements_3          ), //i
    .io_inputs_1_payload_state_elements_4     (poseidonThread_4_io_output_payload_state_elements_4          ), //i
    .io_inputs_1_payload_state_elements_5     (poseidonThread_4_io_output_payload_state_elements_5          ), //i
    .io_inputs_1_payload_state_elements_6     (poseidonThread_4_io_output_payload_state_elements_6          ), //i
    .io_inputs_1_payload_state_elements_7     (poseidonThread_4_io_output_payload_state_elements_7          ), //i
    .io_inputs_1_payload_state_elements_8     (poseidonThread_4_io_output_payload_state_elements_8          ), //i
    .io_inputs_1_payload_state_elements_9     (poseidonThread_4_io_output_payload_state_elements_9          ), //i
    .io_inputs_1_payload_state_elements_10    (poseidonThread_4_io_output_payload_state_elements_10         ), //i
    .io_inputs_1_payload_state_elements_11    (poseidonThread_4_io_output_payload_state_elements_11         ), //i
    .io_inputs_2_valid                        (poseidonThread_5_io_output_valid                             ), //i
    .io_inputs_2_ready                        (DataProcess_matrixAdder_io_inputs_2_ready                    ), //o
    .io_inputs_2_payload_round_index          (poseidonThread_5_io_output_payload_round_index               ), //i
    .io_inputs_2_payload_state_size           (poseidonThread_5_io_output_payload_state_size                ), //i
    .io_inputs_2_payload_state_id             (poseidonThread_5_io_output_payload_state_id                  ), //i
    .io_inputs_2_payload_state_elements_0     (poseidonThread_5_io_output_payload_state_elements_0          ), //i
    .io_inputs_2_payload_state_elements_1     (poseidonThread_5_io_output_payload_state_elements_1          ), //i
    .io_inputs_2_payload_state_elements_2     (poseidonThread_5_io_output_payload_state_elements_2          ), //i
    .io_inputs_2_payload_state_elements_3     (poseidonThread_5_io_output_payload_state_elements_3          ), //i
    .io_inputs_2_payload_state_elements_4     (poseidonThread_5_io_output_payload_state_elements_4          ), //i
    .io_inputs_2_payload_state_elements_5     (poseidonThread_5_io_output_payload_state_elements_5          ), //i
    .io_inputs_2_payload_state_elements_6     (poseidonThread_5_io_output_payload_state_elements_6          ), //i
    .io_inputs_2_payload_state_elements_7     (poseidonThread_5_io_output_payload_state_elements_7          ), //i
    .io_inputs_2_payload_state_elements_8     (poseidonThread_5_io_output_payload_state_elements_8          ), //i
    .io_inputs_2_payload_state_elements_9     (poseidonThread_5_io_output_payload_state_elements_9          ), //i
    .io_inputs_2_payload_state_elements_10    (poseidonThread_5_io_output_payload_state_elements_10         ), //i
    .io_inputs_2_payload_state_elements_11    (poseidonThread_5_io_output_payload_state_elements_11         ), //i
    .io_output_valid                          (DataProcess_matrixAdder_io_output_valid                      ), //o
    .io_output_ready                          (DataProcess_output_ready                                     ), //i
    .io_output_payload_round_index            (DataProcess_matrixAdder_io_output_payload_round_index        ), //o
    .io_output_payload_state_size             (DataProcess_matrixAdder_io_output_payload_state_size         ), //o
    .io_output_payload_state_id               (DataProcess_matrixAdder_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0       (DataProcess_matrixAdder_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1       (DataProcess_matrixAdder_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2       (DataProcess_matrixAdder_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3       (DataProcess_matrixAdder_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4       (DataProcess_matrixAdder_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5       (DataProcess_matrixAdder_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6       (DataProcess_matrixAdder_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7       (DataProcess_matrixAdder_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8       (DataProcess_matrixAdder_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9       (DataProcess_matrixAdder_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10      (DataProcess_matrixAdder_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11      (DataProcess_matrixAdder_io_output_payload_state_elements_11  ), //o
    .clk                                      (clk                                                          ), //i
    .reset                                    (reset                                                        )  //i
  );
  PoseidonThread poseidonThread_3 (
    .io_input_valid                         (DataMux_outputs_0_valid                               ), //i
    .io_input_ready                         (poseidonThread_3_io_input_ready                       ), //o
    .io_input_payload_round_index           (DataMux_outputs_0_payload_round_index                 ), //i
    .io_input_payload_state_index           (DataMux_outputs_0_payload_state_index                 ), //i
    .io_input_payload_state_size            (DataMux_outputs_0_payload_state_size                  ), //i
    .io_input_payload_state_id              (DataMux_outputs_0_payload_state_id                    ), //i
    .io_input_payload_state_element         (DataMux_outputs_0_payload_state_element               ), //i
    .io_output_valid                        (poseidonThread_3_io_output_valid                      ), //o
    .io_output_ready                        (DataProcess_matrixAdder_io_inputs_0_ready             ), //i
    .io_output_payload_round_index          (poseidonThread_3_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (poseidonThread_3_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (poseidonThread_3_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (poseidonThread_3_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (poseidonThread_3_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (poseidonThread_3_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (poseidonThread_3_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (poseidonThread_3_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (poseidonThread_3_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (poseidonThread_3_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (poseidonThread_3_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (poseidonThread_3_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (poseidonThread_3_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (poseidonThread_3_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (poseidonThread_3_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                 ), //i
    .clk                                    (clk                                                   )  //i
  );
  PoseidonThread_1 poseidonThread_4 (
    .io_input_valid                         (DataMux_outputs_1_valid                               ), //i
    .io_input_ready                         (poseidonThread_4_io_input_ready                       ), //o
    .io_input_payload_round_index           (DataMux_outputs_1_payload_round_index                 ), //i
    .io_input_payload_state_index           (DataMux_outputs_1_payload_state_index                 ), //i
    .io_input_payload_state_size            (DataMux_outputs_1_payload_state_size                  ), //i
    .io_input_payload_state_id              (DataMux_outputs_1_payload_state_id                    ), //i
    .io_input_payload_state_element         (DataMux_outputs_1_payload_state_element               ), //i
    .io_output_valid                        (poseidonThread_4_io_output_valid                      ), //o
    .io_output_ready                        (DataProcess_matrixAdder_io_inputs_1_ready             ), //i
    .io_output_payload_round_index          (poseidonThread_4_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (poseidonThread_4_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (poseidonThread_4_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (poseidonThread_4_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (poseidonThread_4_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (poseidonThread_4_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (poseidonThread_4_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (poseidonThread_4_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (poseidonThread_4_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (poseidonThread_4_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (poseidonThread_4_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (poseidonThread_4_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (poseidonThread_4_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (poseidonThread_4_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (poseidonThread_4_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                 ), //i
    .clk                                    (clk                                                   )  //i
  );
  PoseidonThread_2 poseidonThread_5 (
    .io_input_valid                         (DataMux_outputs_2_valid                               ), //i
    .io_input_ready                         (poseidonThread_5_io_input_ready                       ), //o
    .io_input_payload_round_index           (DataMux_outputs_2_payload_round_index                 ), //i
    .io_input_payload_state_index           (DataMux_outputs_2_payload_state_index                 ), //i
    .io_input_payload_state_size            (DataMux_outputs_2_payload_state_size                  ), //i
    .io_input_payload_state_id              (DataMux_outputs_2_payload_state_id                    ), //i
    .io_input_payload_state_element         (DataMux_outputs_2_payload_state_element               ), //i
    .io_output_valid                        (poseidonThread_5_io_output_valid                      ), //o
    .io_output_ready                        (DataProcess_matrixAdder_io_inputs_2_ready             ), //i
    .io_output_payload_round_index          (poseidonThread_5_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (poseidonThread_5_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (poseidonThread_5_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (poseidonThread_5_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (poseidonThread_5_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (poseidonThread_5_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (poseidonThread_5_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (poseidonThread_5_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (poseidonThread_5_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (poseidonThread_5_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (poseidonThread_5_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (poseidonThread_5_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (poseidonThread_5_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (poseidonThread_5_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (poseidonThread_5_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                 ), //i
    .clk                                    (clk                                                   )  //i
  );
  DataLoopbackBuffer loopbackBuffer (
    .io_input_valid                        (DataDeMux_output1_valid                            ), //i
    .io_input_ready                        (loopbackBuffer_io_input_ready                      ), //o
    .io_input_payload_round_index          (DataDeMux_output1_payload_round_index              ), //i
    .io_input_payload_state_size           (DataDeMux_output1_payload_state_size               ), //i
    .io_input_payload_state_id             (DataDeMux_output1_payload_state_id                 ), //i
    .io_input_payload_state_elements_0     (DataDeMux_output1_payload_state_elements_0         ), //i
    .io_input_payload_state_elements_1     (DataDeMux_output1_payload_state_elements_1         ), //i
    .io_input_payload_state_elements_2     (DataDeMux_output1_payload_state_elements_2         ), //i
    .io_input_payload_state_elements_3     (DataDeMux_output1_payload_state_elements_3         ), //i
    .io_input_payload_state_elements_4     (DataDeMux_output1_payload_state_elements_4         ), //i
    .io_input_payload_state_elements_5     (DataDeMux_output1_payload_state_elements_5         ), //i
    .io_input_payload_state_elements_6     (DataDeMux_output1_payload_state_elements_6         ), //i
    .io_input_payload_state_elements_7     (DataDeMux_output1_payload_state_elements_7         ), //i
    .io_input_payload_state_elements_8     (DataDeMux_output1_payload_state_elements_8         ), //i
    .io_input_payload_state_elements_9     (DataDeMux_output1_payload_state_elements_9         ), //i
    .io_input_payload_state_elements_10    (DataDeMux_output1_payload_state_elements_10        ), //i
    .io_input_payload_state_elements_11    (DataDeMux_output1_payload_state_elements_11        ), //i
    .io_outputs_0_valid                    (loopbackBuffer_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (DataMux_inputs0_0_ready                            ), //i
    .io_outputs_0_payload_round_index      (loopbackBuffer_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (loopbackBuffer_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (loopbackBuffer_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (loopbackBuffer_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (loopbackBuffer_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (loopbackBuffer_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (DataMux_inputs0_1_ready                            ), //i
    .io_outputs_1_payload_round_index      (loopbackBuffer_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (loopbackBuffer_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (loopbackBuffer_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (loopbackBuffer_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (loopbackBuffer_io_outputs_1_payload_state_element  ), //o
    .io_outputs_2_valid                    (loopbackBuffer_io_outputs_2_valid                  ), //o
    .io_outputs_2_ready                    (DataMux_inputs0_2_ready                            ), //i
    .io_outputs_2_payload_round_index      (loopbackBuffer_io_outputs_2_payload_round_index    ), //o
    .io_outputs_2_payload_state_index      (loopbackBuffer_io_outputs_2_payload_state_index    ), //o
    .io_outputs_2_payload_state_size       (loopbackBuffer_io_outputs_2_payload_state_size     ), //o
    .io_outputs_2_payload_state_id         (loopbackBuffer_io_outputs_2_payload_state_id       ), //o
    .io_outputs_2_payload_state_element    (loopbackBuffer_io_outputs_2_payload_state_element  ), //o
    .io_residue                            (loopbackBuffer_io_residue                          ), //o
    .clk                                   (clk                                                ), //i
    .reset                                 (reset                                              )  //i
  );
  AXI4StreamTransmitter transmitter (
    .io_input_valid                    (DataDeMux_output0_valid                  ), //i
    .io_input_ready                    (transmitter_io_input_ready               ), //o
    .io_input_payload_state_id         (DataDeMux_output0_payload_state_id       ), //i
    .io_input_payload_state_element    (DataDeMux_output0_payload_state_element  ), //i
    .io_output_valid                   (transmitter_io_output_valid              ), //o
    .io_output_ready                   (io_output_ready                          ), //i
    .io_output_last                    (transmitter_io_output_last               ), //o
    .io_output_payload                 (transmitter_io_output_payload            ), //o
    .clk                               (clk                                      ), //i
    .reset                             (reset                                    )  //i
  );
  assign io_input_ready = receiver_io_input_ready;
  assign receiver_io_outputs_0_ready = (! receiver_io_outputs_0_rValid);
  assign receiver_io_outputs_0_s2mPipe_valid = (receiver_io_outputs_0_valid || receiver_io_outputs_0_rValid);
  assign receiver_io_outputs_0_s2mPipe_payload_round_index = (receiver_io_outputs_0_rValid ? receiver_io_outputs_0_rData_round_index : receiver_io_outputs_0_payload_round_index);
  assign receiver_io_outputs_0_s2mPipe_payload_state_index = (receiver_io_outputs_0_rValid ? receiver_io_outputs_0_rData_state_index : receiver_io_outputs_0_payload_state_index);
  assign receiver_io_outputs_0_s2mPipe_payload_state_size = (receiver_io_outputs_0_rValid ? receiver_io_outputs_0_rData_state_size : receiver_io_outputs_0_payload_state_size);
  assign receiver_io_outputs_0_s2mPipe_payload_state_id = (receiver_io_outputs_0_rValid ? receiver_io_outputs_0_rData_state_id : receiver_io_outputs_0_payload_state_id);
  assign receiver_io_outputs_0_s2mPipe_payload_state_element = (receiver_io_outputs_0_rValid ? receiver_io_outputs_0_rData_state_element : receiver_io_outputs_0_payload_state_element);
  always @(*) begin
    receiver_io_outputs_0_s2mPipe_ready = receiver_io_outputs_0_s2mPipe_m2sPipe_ready;
    if(when_Stream_l342) begin
      receiver_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! receiver_io_outputs_0_s2mPipe_m2sPipe_valid);
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_valid = receiver_io_outputs_0_s2mPipe_rValid;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_payload_round_index = receiver_io_outputs_0_s2mPipe_rData_round_index;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_index = receiver_io_outputs_0_s2mPipe_rData_state_index;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_size = receiver_io_outputs_0_s2mPipe_rData_state_size;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_id = receiver_io_outputs_0_s2mPipe_rData_state_id;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_element = receiver_io_outputs_0_s2mPipe_rData_state_element;
  assign DataMux_inputs1_temp_0_valid = receiver_io_outputs_0_s2mPipe_m2sPipe_valid;
  assign receiver_io_outputs_0_s2mPipe_m2sPipe_ready = DataMux_inputs1_temp_0_ready;
  assign DataMux_inputs1_temp_0_payload_round_index = receiver_io_outputs_0_s2mPipe_m2sPipe_payload_round_index;
  assign DataMux_inputs1_temp_0_payload_state_index = receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_index;
  assign DataMux_inputs1_temp_0_payload_state_size = receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_size;
  assign DataMux_inputs1_temp_0_payload_state_id = receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_id;
  assign DataMux_inputs1_temp_0_payload_state_element = receiver_io_outputs_0_s2mPipe_m2sPipe_payload_state_element;
  assign receiver_io_outputs_1_ready = (! receiver_io_outputs_1_rValid);
  assign receiver_io_outputs_1_s2mPipe_valid = (receiver_io_outputs_1_valid || receiver_io_outputs_1_rValid);
  assign receiver_io_outputs_1_s2mPipe_payload_round_index = (receiver_io_outputs_1_rValid ? receiver_io_outputs_1_rData_round_index : receiver_io_outputs_1_payload_round_index);
  assign receiver_io_outputs_1_s2mPipe_payload_state_index = (receiver_io_outputs_1_rValid ? receiver_io_outputs_1_rData_state_index : receiver_io_outputs_1_payload_state_index);
  assign receiver_io_outputs_1_s2mPipe_payload_state_size = (receiver_io_outputs_1_rValid ? receiver_io_outputs_1_rData_state_size : receiver_io_outputs_1_payload_state_size);
  assign receiver_io_outputs_1_s2mPipe_payload_state_id = (receiver_io_outputs_1_rValid ? receiver_io_outputs_1_rData_state_id : receiver_io_outputs_1_payload_state_id);
  assign receiver_io_outputs_1_s2mPipe_payload_state_element = (receiver_io_outputs_1_rValid ? receiver_io_outputs_1_rData_state_element : receiver_io_outputs_1_payload_state_element);
  always @(*) begin
    receiver_io_outputs_1_s2mPipe_ready = receiver_io_outputs_1_s2mPipe_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      receiver_io_outputs_1_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! receiver_io_outputs_1_s2mPipe_m2sPipe_valid);
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_valid = receiver_io_outputs_1_s2mPipe_rValid;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_payload_round_index = receiver_io_outputs_1_s2mPipe_rData_round_index;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_index = receiver_io_outputs_1_s2mPipe_rData_state_index;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_size = receiver_io_outputs_1_s2mPipe_rData_state_size;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_id = receiver_io_outputs_1_s2mPipe_rData_state_id;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_element = receiver_io_outputs_1_s2mPipe_rData_state_element;
  assign DataMux_inputs1_temp_1_valid = receiver_io_outputs_1_s2mPipe_m2sPipe_valid;
  assign receiver_io_outputs_1_s2mPipe_m2sPipe_ready = DataMux_inputs1_temp_1_ready;
  assign DataMux_inputs1_temp_1_payload_round_index = receiver_io_outputs_1_s2mPipe_m2sPipe_payload_round_index;
  assign DataMux_inputs1_temp_1_payload_state_index = receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_index;
  assign DataMux_inputs1_temp_1_payload_state_size = receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_size;
  assign DataMux_inputs1_temp_1_payload_state_id = receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_id;
  assign DataMux_inputs1_temp_1_payload_state_element = receiver_io_outputs_1_s2mPipe_m2sPipe_payload_state_element;
  assign receiver_io_outputs_2_ready = (! receiver_io_outputs_2_rValid);
  assign receiver_io_outputs_2_s2mPipe_valid = (receiver_io_outputs_2_valid || receiver_io_outputs_2_rValid);
  assign receiver_io_outputs_2_s2mPipe_payload_round_index = (receiver_io_outputs_2_rValid ? receiver_io_outputs_2_rData_round_index : receiver_io_outputs_2_payload_round_index);
  assign receiver_io_outputs_2_s2mPipe_payload_state_index = (receiver_io_outputs_2_rValid ? receiver_io_outputs_2_rData_state_index : receiver_io_outputs_2_payload_state_index);
  assign receiver_io_outputs_2_s2mPipe_payload_state_size = (receiver_io_outputs_2_rValid ? receiver_io_outputs_2_rData_state_size : receiver_io_outputs_2_payload_state_size);
  assign receiver_io_outputs_2_s2mPipe_payload_state_id = (receiver_io_outputs_2_rValid ? receiver_io_outputs_2_rData_state_id : receiver_io_outputs_2_payload_state_id);
  assign receiver_io_outputs_2_s2mPipe_payload_state_element = (receiver_io_outputs_2_rValid ? receiver_io_outputs_2_rData_state_element : receiver_io_outputs_2_payload_state_element);
  always @(*) begin
    receiver_io_outputs_2_s2mPipe_ready = receiver_io_outputs_2_s2mPipe_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      receiver_io_outputs_2_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! receiver_io_outputs_2_s2mPipe_m2sPipe_valid);
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_valid = receiver_io_outputs_2_s2mPipe_rValid;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_payload_round_index = receiver_io_outputs_2_s2mPipe_rData_round_index;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_index = receiver_io_outputs_2_s2mPipe_rData_state_index;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_size = receiver_io_outputs_2_s2mPipe_rData_state_size;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_id = receiver_io_outputs_2_s2mPipe_rData_state_id;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_element = receiver_io_outputs_2_s2mPipe_rData_state_element;
  assign DataMux_inputs1_temp_2_valid = receiver_io_outputs_2_s2mPipe_m2sPipe_valid;
  assign receiver_io_outputs_2_s2mPipe_m2sPipe_ready = DataMux_inputs1_temp_2_ready;
  assign DataMux_inputs1_temp_2_payload_round_index = receiver_io_outputs_2_s2mPipe_m2sPipe_payload_round_index;
  assign DataMux_inputs1_temp_2_payload_state_index = receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_index;
  assign DataMux_inputs1_temp_2_payload_state_size = receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_size;
  assign DataMux_inputs1_temp_2_payload_state_id = receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_id;
  assign DataMux_inputs1_temp_2_payload_state_element = receiver_io_outputs_2_s2mPipe_m2sPipe_payload_state_element;
  assign _zz_DataMux_inputs1_temp_0_ready = (_zz__zz_DataMux_inputs1_temp_0_ready <= DataMux_residue);
  assign DataMux_inputs1_0_valid = (DataMux_inputs1_temp_0_valid && _zz_DataMux_inputs1_temp_0_ready);
  assign DataMux_inputs1_temp_0_ready = (DataMux_inputs1_0_ready && _zz_DataMux_inputs1_temp_0_ready);
  assign DataMux_inputs1_0_payload_round_index = DataMux_inputs1_temp_0_payload_round_index;
  assign DataMux_inputs1_0_payload_state_index = DataMux_inputs1_temp_0_payload_state_index;
  assign DataMux_inputs1_0_payload_state_size = DataMux_inputs1_temp_0_payload_state_size;
  assign DataMux_inputs1_0_payload_state_id = DataMux_inputs1_temp_0_payload_state_id;
  assign DataMux_inputs1_0_payload_state_element = DataMux_inputs1_temp_0_payload_state_element;
  assign _zz_DataMux_inputs1_temp_1_ready = (_zz__zz_DataMux_inputs1_temp_1_ready <= DataMux_residue);
  assign DataMux_inputs1_1_valid = (DataMux_inputs1_temp_1_valid && _zz_DataMux_inputs1_temp_1_ready);
  assign DataMux_inputs1_temp_1_ready = (DataMux_inputs1_1_ready && _zz_DataMux_inputs1_temp_1_ready);
  assign DataMux_inputs1_1_payload_round_index = DataMux_inputs1_temp_1_payload_round_index;
  assign DataMux_inputs1_1_payload_state_index = DataMux_inputs1_temp_1_payload_state_index;
  assign DataMux_inputs1_1_payload_state_size = DataMux_inputs1_temp_1_payload_state_size;
  assign DataMux_inputs1_1_payload_state_id = DataMux_inputs1_temp_1_payload_state_id;
  assign DataMux_inputs1_1_payload_state_element = DataMux_inputs1_temp_1_payload_state_element;
  assign _zz_DataMux_inputs1_temp_2_ready = (_zz__zz_DataMux_inputs1_temp_2_ready <= DataMux_residue);
  assign DataMux_inputs1_2_valid = (DataMux_inputs1_temp_2_valid && _zz_DataMux_inputs1_temp_2_ready);
  assign DataMux_inputs1_temp_2_ready = (DataMux_inputs1_2_ready && _zz_DataMux_inputs1_temp_2_ready);
  assign DataMux_inputs1_2_payload_round_index = DataMux_inputs1_temp_2_payload_round_index;
  assign DataMux_inputs1_2_payload_state_index = DataMux_inputs1_temp_2_payload_state_index;
  assign DataMux_inputs1_2_payload_state_size = DataMux_inputs1_temp_2_payload_state_size;
  assign DataMux_inputs1_2_payload_state_id = DataMux_inputs1_temp_2_payload_state_id;
  assign DataMux_inputs1_2_payload_state_element = DataMux_inputs1_temp_2_payload_state_element;
  assign DataMux_inputs0_0_ready = streamArbiter_12_io_inputs_0_ready;
  assign DataMux_inputs1_0_ready = streamArbiter_12_io_inputs_1_ready;
  assign DataMux_outputs_0_valid = streamArbiter_12_io_output_valid;
  assign DataMux_outputs_0_payload_round_index = streamArbiter_12_io_output_payload_round_index;
  assign DataMux_outputs_0_payload_state_index = streamArbiter_12_io_output_payload_state_index;
  assign DataMux_outputs_0_payload_state_size = streamArbiter_12_io_output_payload_state_size;
  assign DataMux_outputs_0_payload_state_id = streamArbiter_12_io_output_payload_state_id;
  assign DataMux_outputs_0_payload_state_element = streamArbiter_12_io_output_payload_state_element;
  assign DataMux_inputs0_1_ready = streamArbiter_13_io_inputs_0_ready;
  assign DataMux_inputs1_1_ready = streamArbiter_13_io_inputs_1_ready;
  assign DataMux_outputs_1_valid = streamArbiter_13_io_output_valid;
  assign DataMux_outputs_1_payload_round_index = streamArbiter_13_io_output_payload_round_index;
  assign DataMux_outputs_1_payload_state_index = streamArbiter_13_io_output_payload_state_index;
  assign DataMux_outputs_1_payload_state_size = streamArbiter_13_io_output_payload_state_size;
  assign DataMux_outputs_1_payload_state_id = streamArbiter_13_io_output_payload_state_id;
  assign DataMux_outputs_1_payload_state_element = streamArbiter_13_io_output_payload_state_element;
  assign DataMux_inputs0_2_ready = streamArbiter_14_io_inputs_0_ready;
  assign DataMux_inputs1_2_ready = streamArbiter_14_io_inputs_1_ready;
  assign DataMux_outputs_2_valid = streamArbiter_14_io_output_valid;
  assign DataMux_outputs_2_payload_round_index = streamArbiter_14_io_output_payload_round_index;
  assign DataMux_outputs_2_payload_state_index = streamArbiter_14_io_output_payload_state_index;
  assign DataMux_outputs_2_payload_state_size = streamArbiter_14_io_output_payload_state_size;
  assign DataMux_outputs_2_payload_state_id = streamArbiter_14_io_output_payload_state_id;
  assign DataMux_outputs_2_payload_state_element = streamArbiter_14_io_output_payload_state_element;
  assign DataProcess_output_valid = DataProcess_matrixAdder_io_output_valid;
  assign DataProcess_output_payload_round_index = DataProcess_matrixAdder_io_output_payload_round_index;
  assign DataProcess_output_payload_state_size = DataProcess_matrixAdder_io_output_payload_state_size;
  assign DataProcess_output_payload_state_id = DataProcess_matrixAdder_io_output_payload_state_id;
  assign DataProcess_output_payload_state_elements_0 = DataProcess_matrixAdder_io_output_payload_state_elements_0;
  assign DataProcess_output_payload_state_elements_1 = DataProcess_matrixAdder_io_output_payload_state_elements_1;
  assign DataProcess_output_payload_state_elements_2 = DataProcess_matrixAdder_io_output_payload_state_elements_2;
  assign DataProcess_output_payload_state_elements_3 = DataProcess_matrixAdder_io_output_payload_state_elements_3;
  assign DataProcess_output_payload_state_elements_4 = DataProcess_matrixAdder_io_output_payload_state_elements_4;
  assign DataProcess_output_payload_state_elements_5 = DataProcess_matrixAdder_io_output_payload_state_elements_5;
  assign DataProcess_output_payload_state_elements_6 = DataProcess_matrixAdder_io_output_payload_state_elements_6;
  assign DataProcess_output_payload_state_elements_7 = DataProcess_matrixAdder_io_output_payload_state_elements_7;
  assign DataProcess_output_payload_state_elements_8 = DataProcess_matrixAdder_io_output_payload_state_elements_8;
  assign DataProcess_output_payload_state_elements_9 = DataProcess_matrixAdder_io_output_payload_state_elements_9;
  assign DataProcess_output_payload_state_elements_10 = DataProcess_matrixAdder_io_output_payload_state_elements_10;
  assign DataProcess_output_payload_state_elements_11 = DataProcess_matrixAdder_io_output_payload_state_elements_11;
  assign DataMux_outputs_0_ready = poseidonThread_3_io_input_ready;
  assign DataMux_outputs_1_ready = poseidonThread_4_io_input_ready;
  assign DataMux_outputs_2_ready = poseidonThread_5_io_input_ready;
  assign DataDeMux_output0_valid = (DataProcess_output_valid && DataDeMux_select[0]);
  assign DataDeMux_output1_valid = (DataProcess_output_valid && DataDeMux_select[1]);
  assign DataProcess_output_ready = ((DataDeMux_output0_ready && DataDeMux_select[0]) || (DataDeMux_output1_ready && DataDeMux_select[1]));
  assign DataDeMux_output0_payload_state_id = DataProcess_output_payload_state_id;
  assign DataDeMux_output0_payload_state_element = DataProcess_output_payload_state_elements_1;
  always @(*) begin
    DataDeMux_output1_payload_round_index = DataProcess_output_payload_round_index;
    DataDeMux_output1_payload_round_index = (DataProcess_output_payload_round_index + 7'h01);
  end

  assign DataDeMux_output1_payload_state_size = DataProcess_output_payload_state_size;
  assign DataDeMux_output1_payload_state_id = DataProcess_output_payload_state_id;
  assign DataDeMux_output1_payload_state_elements_0 = DataProcess_output_payload_state_elements_0;
  assign DataDeMux_output1_payload_state_elements_1 = DataProcess_output_payload_state_elements_1;
  assign DataDeMux_output1_payload_state_elements_2 = DataProcess_output_payload_state_elements_2;
  assign DataDeMux_output1_payload_state_elements_3 = DataProcess_output_payload_state_elements_3;
  assign DataDeMux_output1_payload_state_elements_4 = DataProcess_output_payload_state_elements_4;
  assign DataDeMux_output1_payload_state_elements_5 = DataProcess_output_payload_state_elements_5;
  assign DataDeMux_output1_payload_state_elements_6 = DataProcess_output_payload_state_elements_6;
  assign DataDeMux_output1_payload_state_elements_7 = DataProcess_output_payload_state_elements_7;
  assign DataDeMux_output1_payload_state_elements_8 = DataProcess_output_payload_state_elements_8;
  assign DataDeMux_output1_payload_state_elements_9 = DataProcess_output_payload_state_elements_9;
  assign DataDeMux_output1_payload_state_elements_10 = DataProcess_output_payload_state_elements_10;
  assign DataDeMux_output1_payload_state_elements_11 = DataProcess_output_payload_state_elements_11;
  always @(*) begin
    case(DataProcess_output_payload_state_size)
      4'b0011 : begin
        DataDeMux_select[0] = (DataProcess_output_payload_round_index == 7'h3e);
        DataDeMux_select[1] = (DataProcess_output_payload_round_index < 7'h3e);
      end
      4'b0101 : begin
        DataDeMux_select[0] = (DataProcess_output_payload_round_index == 7'h3f);
        DataDeMux_select[1] = (DataProcess_output_payload_round_index < 7'h3f);
      end
      4'b1001 : begin
        DataDeMux_select[0] = (DataProcess_output_payload_round_index == 7'h40);
        DataDeMux_select[1] = (DataProcess_output_payload_round_index < 7'h40);
      end
      4'b1100 : begin
        DataDeMux_select[0] = (DataProcess_output_payload_round_index == 7'h40);
        DataDeMux_select[1] = (DataProcess_output_payload_round_index < 7'h40);
      end
      default : begin
        DataDeMux_select = 2'b00;
      end
    endcase
  end

  assign DataDeMux_output1_ready = loopbackBuffer_io_input_ready;
  assign DataMux_inputs0_0_valid = loopbackBuffer_io_outputs_0_valid;
  assign DataMux_inputs0_0_payload_round_index = loopbackBuffer_io_outputs_0_payload_round_index;
  assign DataMux_inputs0_0_payload_state_index = loopbackBuffer_io_outputs_0_payload_state_index;
  assign DataMux_inputs0_0_payload_state_size = loopbackBuffer_io_outputs_0_payload_state_size;
  assign DataMux_inputs0_0_payload_state_id = loopbackBuffer_io_outputs_0_payload_state_id;
  assign DataMux_inputs0_0_payload_state_element = loopbackBuffer_io_outputs_0_payload_state_element;
  assign DataMux_inputs0_1_valid = loopbackBuffer_io_outputs_1_valid;
  assign DataMux_inputs0_1_payload_round_index = loopbackBuffer_io_outputs_1_payload_round_index;
  assign DataMux_inputs0_1_payload_state_index = loopbackBuffer_io_outputs_1_payload_state_index;
  assign DataMux_inputs0_1_payload_state_size = loopbackBuffer_io_outputs_1_payload_state_size;
  assign DataMux_inputs0_1_payload_state_id = loopbackBuffer_io_outputs_1_payload_state_id;
  assign DataMux_inputs0_1_payload_state_element = loopbackBuffer_io_outputs_1_payload_state_element;
  assign DataMux_inputs0_2_valid = loopbackBuffer_io_outputs_2_valid;
  assign DataMux_inputs0_2_payload_round_index = loopbackBuffer_io_outputs_2_payload_round_index;
  assign DataMux_inputs0_2_payload_state_index = loopbackBuffer_io_outputs_2_payload_state_index;
  assign DataMux_inputs0_2_payload_state_size = loopbackBuffer_io_outputs_2_payload_state_size;
  assign DataMux_inputs0_2_payload_state_id = loopbackBuffer_io_outputs_2_payload_state_id;
  assign DataMux_inputs0_2_payload_state_element = loopbackBuffer_io_outputs_2_payload_state_element;
  assign DataMux_residue = loopbackBuffer_io_residue;
  assign DataDeMux_output0_ready = transmitter_io_input_ready;
  assign io_output_valid = transmitter_io_output_valid;
  assign io_output_last = transmitter_io_output_last;
  assign io_output_payload = transmitter_io_output_payload;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      receiver_io_outputs_0_rValid <= 1'b0;
      receiver_io_outputs_0_s2mPipe_rValid <= 1'b0;
      receiver_io_outputs_1_rValid <= 1'b0;
      receiver_io_outputs_1_s2mPipe_rValid <= 1'b0;
      receiver_io_outputs_2_rValid <= 1'b0;
      receiver_io_outputs_2_s2mPipe_rValid <= 1'b0;
    end else begin
      if(receiver_io_outputs_0_valid) begin
        receiver_io_outputs_0_rValid <= 1'b1;
      end
      if(receiver_io_outputs_0_s2mPipe_ready) begin
        receiver_io_outputs_0_rValid <= 1'b0;
      end
      if(receiver_io_outputs_0_s2mPipe_ready) begin
        receiver_io_outputs_0_s2mPipe_rValid <= receiver_io_outputs_0_s2mPipe_valid;
      end
      if(receiver_io_outputs_1_valid) begin
        receiver_io_outputs_1_rValid <= 1'b1;
      end
      if(receiver_io_outputs_1_s2mPipe_ready) begin
        receiver_io_outputs_1_rValid <= 1'b0;
      end
      if(receiver_io_outputs_1_s2mPipe_ready) begin
        receiver_io_outputs_1_s2mPipe_rValid <= receiver_io_outputs_1_s2mPipe_valid;
      end
      if(receiver_io_outputs_2_valid) begin
        receiver_io_outputs_2_rValid <= 1'b1;
      end
      if(receiver_io_outputs_2_s2mPipe_ready) begin
        receiver_io_outputs_2_rValid <= 1'b0;
      end
      if(receiver_io_outputs_2_s2mPipe_ready) begin
        receiver_io_outputs_2_s2mPipe_rValid <= receiver_io_outputs_2_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(receiver_io_outputs_0_ready) begin
      receiver_io_outputs_0_rData_round_index <= receiver_io_outputs_0_payload_round_index;
      receiver_io_outputs_0_rData_state_index <= receiver_io_outputs_0_payload_state_index;
      receiver_io_outputs_0_rData_state_size <= receiver_io_outputs_0_payload_state_size;
      receiver_io_outputs_0_rData_state_id <= receiver_io_outputs_0_payload_state_id;
      receiver_io_outputs_0_rData_state_element <= receiver_io_outputs_0_payload_state_element;
    end
    if(receiver_io_outputs_0_s2mPipe_ready) begin
      receiver_io_outputs_0_s2mPipe_rData_round_index <= receiver_io_outputs_0_s2mPipe_payload_round_index;
      receiver_io_outputs_0_s2mPipe_rData_state_index <= receiver_io_outputs_0_s2mPipe_payload_state_index;
      receiver_io_outputs_0_s2mPipe_rData_state_size <= receiver_io_outputs_0_s2mPipe_payload_state_size;
      receiver_io_outputs_0_s2mPipe_rData_state_id <= receiver_io_outputs_0_s2mPipe_payload_state_id;
      receiver_io_outputs_0_s2mPipe_rData_state_element <= receiver_io_outputs_0_s2mPipe_payload_state_element;
    end
    if(receiver_io_outputs_1_ready) begin
      receiver_io_outputs_1_rData_round_index <= receiver_io_outputs_1_payload_round_index;
      receiver_io_outputs_1_rData_state_index <= receiver_io_outputs_1_payload_state_index;
      receiver_io_outputs_1_rData_state_size <= receiver_io_outputs_1_payload_state_size;
      receiver_io_outputs_1_rData_state_id <= receiver_io_outputs_1_payload_state_id;
      receiver_io_outputs_1_rData_state_element <= receiver_io_outputs_1_payload_state_element;
    end
    if(receiver_io_outputs_1_s2mPipe_ready) begin
      receiver_io_outputs_1_s2mPipe_rData_round_index <= receiver_io_outputs_1_s2mPipe_payload_round_index;
      receiver_io_outputs_1_s2mPipe_rData_state_index <= receiver_io_outputs_1_s2mPipe_payload_state_index;
      receiver_io_outputs_1_s2mPipe_rData_state_size <= receiver_io_outputs_1_s2mPipe_payload_state_size;
      receiver_io_outputs_1_s2mPipe_rData_state_id <= receiver_io_outputs_1_s2mPipe_payload_state_id;
      receiver_io_outputs_1_s2mPipe_rData_state_element <= receiver_io_outputs_1_s2mPipe_payload_state_element;
    end
    if(receiver_io_outputs_2_ready) begin
      receiver_io_outputs_2_rData_round_index <= receiver_io_outputs_2_payload_round_index;
      receiver_io_outputs_2_rData_state_index <= receiver_io_outputs_2_payload_state_index;
      receiver_io_outputs_2_rData_state_size <= receiver_io_outputs_2_payload_state_size;
      receiver_io_outputs_2_rData_state_id <= receiver_io_outputs_2_payload_state_id;
      receiver_io_outputs_2_rData_state_element <= receiver_io_outputs_2_payload_state_element;
    end
    if(receiver_io_outputs_2_s2mPipe_ready) begin
      receiver_io_outputs_2_s2mPipe_rData_round_index <= receiver_io_outputs_2_s2mPipe_payload_round_index;
      receiver_io_outputs_2_s2mPipe_rData_state_index <= receiver_io_outputs_2_s2mPipe_payload_state_index;
      receiver_io_outputs_2_s2mPipe_rData_state_size <= receiver_io_outputs_2_s2mPipe_payload_state_size;
      receiver_io_outputs_2_s2mPipe_rData_state_id <= receiver_io_outputs_2_s2mPipe_payload_state_id;
      receiver_io_outputs_2_s2mPipe_rData_state_element <= receiver_io_outputs_2_s2mPipe_payload_state_element;
    end
  end


endmodule

module AXI4StreamTransmitter (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_last,
  output     [254:0]  io_output_payload,
  input               clk,
  input               reset
);
  wire                streamMux_7_io_output_ready;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_0_payload_state_element;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_outputs_2_valid;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_2_payload_state_element;
  wire                streamDemux_7_io_outputs_3_valid;
  wire       [6:0]    streamDemux_7_io_outputs_3_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_3_payload_state_element;
  wire                streamDemux_7_io_outputs_4_valid;
  wire       [6:0]    streamDemux_7_io_outputs_4_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_4_payload_state_element;
  wire                streamDemux_7_io_outputs_5_valid;
  wire       [6:0]    streamDemux_7_io_outputs_5_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_5_payload_state_element;
  wire                streamMux_7_io_inputs_0_ready;
  wire                streamMux_7_io_inputs_1_ready;
  wire                streamMux_7_io_inputs_2_ready;
  wire                streamMux_7_io_inputs_3_ready;
  wire                streamMux_7_io_inputs_4_ready;
  wire                streamMux_7_io_inputs_5_ready;
  wire                streamMux_7_io_output_valid;
  wire       [6:0]    streamMux_7_io_output_payload_state_id;
  wire       [254:0]  streamMux_7_io_output_payload_state_element;
  wire       [5:0]    _zz__zz_demux_select_1;
  reg        [6:0]    idCounter;
  wire                when_AXI4StreamInterface_l211;
  wire                input_demux_0_valid;
  reg                 input_demux_0_ready;
  wire       [6:0]    input_demux_0_payload_state_id;
  wire       [254:0]  input_demux_0_payload_state_element;
  wire                input_demux_1_valid;
  reg                 input_demux_1_ready;
  wire       [6:0]    input_demux_1_payload_state_id;
  wire       [254:0]  input_demux_1_payload_state_element;
  wire                input_demux_2_valid;
  reg                 input_demux_2_ready;
  wire       [6:0]    input_demux_2_payload_state_id;
  wire       [254:0]  input_demux_2_payload_state_element;
  wire                input_demux_3_valid;
  reg                 input_demux_3_ready;
  wire       [6:0]    input_demux_3_payload_state_id;
  wire       [254:0]  input_demux_3_payload_state_element;
  wire                input_demux_4_valid;
  reg                 input_demux_4_ready;
  wire       [6:0]    input_demux_4_payload_state_id;
  wire       [254:0]  input_demux_4_payload_state_element;
  wire                input_demux_5_valid;
  reg                 input_demux_5_ready;
  wire       [6:0]    input_demux_5_payload_state_id;
  wire       [254:0]  input_demux_5_payload_state_element;
  wire       [5:0]    _zz_demux_select;
  wire       [5:0]    _zz_demux_select_1;
  wire                _zz_demux_select_2;
  wire                _zz_demux_select_3;
  wire                _zz_demux_select_4;
  wire                _zz_demux_select_5;
  wire                _zz_demux_select_6;
  wire       [2:0]    demux_select;
  wire                buffer_0_valid;
  wire                buffer_0_ready;
  wire       [6:0]    buffer_0_payload_state_id;
  wire       [254:0]  buffer_0_payload_state_element;
  reg                 input_demux_0_rValid;
  reg        [6:0]    input_demux_0_rData_state_id;
  reg        [254:0]  input_demux_0_rData_state_element;
  wire                when_Stream_l342;
  wire                buffer_1_valid;
  wire                buffer_1_ready;
  wire       [6:0]    buffer_1_payload_state_id;
  wire       [254:0]  buffer_1_payload_state_element;
  reg                 input_demux_1_rValid;
  reg        [6:0]    input_demux_1_rData_state_id;
  reg        [254:0]  input_demux_1_rData_state_element;
  wire                when_Stream_l342_1;
  wire                buffer_2_valid;
  wire                buffer_2_ready;
  wire       [6:0]    buffer_2_payload_state_id;
  wire       [254:0]  buffer_2_payload_state_element;
  reg                 input_demux_2_rValid;
  reg        [6:0]    input_demux_2_rData_state_id;
  reg        [254:0]  input_demux_2_rData_state_element;
  wire                when_Stream_l342_2;
  wire                buffer_3_valid;
  wire                buffer_3_ready;
  wire       [6:0]    buffer_3_payload_state_id;
  wire       [254:0]  buffer_3_payload_state_element;
  reg                 input_demux_3_rValid;
  reg        [6:0]    input_demux_3_rData_state_id;
  reg        [254:0]  input_demux_3_rData_state_element;
  wire                when_Stream_l342_3;
  wire                buffer_4_valid;
  wire                buffer_4_ready;
  wire       [6:0]    buffer_4_payload_state_id;
  wire       [254:0]  buffer_4_payload_state_element;
  reg                 input_demux_4_rValid;
  reg        [6:0]    input_demux_4_rData_state_id;
  reg        [254:0]  input_demux_4_rData_state_element;
  wire                when_Stream_l342_4;
  wire                buffer_5_valid;
  wire                buffer_5_ready;
  wire       [6:0]    buffer_5_payload_state_id;
  wire       [254:0]  buffer_5_payload_state_element;
  reg                 input_demux_5_rValid;
  reg        [6:0]    input_demux_5_rData_state_id;
  reg        [254:0]  input_demux_5_rData_state_element;
  wire                when_Stream_l342_5;
  wire                _zz_select;
  wire                _zz_select_1;
  wire                _zz_select_2;
  wire                _zz_select_3;
  wire                _zz_select_4;
  wire       [2:0]    select_1;

  assign _zz__zz_demux_select_1 = (_zz_demux_select - 6'h01);
  StreamDemux_6 streamDemux_7 (
    .io_select                             (demux_select                                      ), //i
    .io_input_valid                        (io_input_valid                                    ), //i
    .io_input_ready                        (streamDemux_7_io_input_ready                      ), //o
    .io_input_payload_state_id             (io_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (io_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (streamDemux_7_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (input_demux_0_ready                               ), //i
    .io_outputs_0_payload_state_id         (streamDemux_7_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (streamDemux_7_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (streamDemux_7_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (input_demux_1_ready                               ), //i
    .io_outputs_1_payload_state_id         (streamDemux_7_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (streamDemux_7_io_outputs_1_payload_state_element  ), //o
    .io_outputs_2_valid                    (streamDemux_7_io_outputs_2_valid                  ), //o
    .io_outputs_2_ready                    (input_demux_2_ready                               ), //i
    .io_outputs_2_payload_state_id         (streamDemux_7_io_outputs_2_payload_state_id       ), //o
    .io_outputs_2_payload_state_element    (streamDemux_7_io_outputs_2_payload_state_element  ), //o
    .io_outputs_3_valid                    (streamDemux_7_io_outputs_3_valid                  ), //o
    .io_outputs_3_ready                    (input_demux_3_ready                               ), //i
    .io_outputs_3_payload_state_id         (streamDemux_7_io_outputs_3_payload_state_id       ), //o
    .io_outputs_3_payload_state_element    (streamDemux_7_io_outputs_3_payload_state_element  ), //o
    .io_outputs_4_valid                    (streamDemux_7_io_outputs_4_valid                  ), //o
    .io_outputs_4_ready                    (input_demux_4_ready                               ), //i
    .io_outputs_4_payload_state_id         (streamDemux_7_io_outputs_4_payload_state_id       ), //o
    .io_outputs_4_payload_state_element    (streamDemux_7_io_outputs_4_payload_state_element  ), //o
    .io_outputs_5_valid                    (streamDemux_7_io_outputs_5_valid                  ), //o
    .io_outputs_5_ready                    (input_demux_5_ready                               ), //i
    .io_outputs_5_payload_state_id         (streamDemux_7_io_outputs_5_payload_state_id       ), //o
    .io_outputs_5_payload_state_element    (streamDemux_7_io_outputs_5_payload_state_element  )  //o
  );
  StreamMux_6 streamMux_7 (
    .io_select                            (select_1                                     ), //i
    .io_inputs_0_valid                    (buffer_0_valid                               ), //i
    .io_inputs_0_ready                    (streamMux_7_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_state_id         (buffer_0_payload_state_id                    ), //i
    .io_inputs_0_payload_state_element    (buffer_0_payload_state_element               ), //i
    .io_inputs_1_valid                    (buffer_1_valid                               ), //i
    .io_inputs_1_ready                    (streamMux_7_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_state_id         (buffer_1_payload_state_id                    ), //i
    .io_inputs_1_payload_state_element    (buffer_1_payload_state_element               ), //i
    .io_inputs_2_valid                    (buffer_2_valid                               ), //i
    .io_inputs_2_ready                    (streamMux_7_io_inputs_2_ready                ), //o
    .io_inputs_2_payload_state_id         (buffer_2_payload_state_id                    ), //i
    .io_inputs_2_payload_state_element    (buffer_2_payload_state_element               ), //i
    .io_inputs_3_valid                    (buffer_3_valid                               ), //i
    .io_inputs_3_ready                    (streamMux_7_io_inputs_3_ready                ), //o
    .io_inputs_3_payload_state_id         (buffer_3_payload_state_id                    ), //i
    .io_inputs_3_payload_state_element    (buffer_3_payload_state_element               ), //i
    .io_inputs_4_valid                    (buffer_4_valid                               ), //i
    .io_inputs_4_ready                    (streamMux_7_io_inputs_4_ready                ), //o
    .io_inputs_4_payload_state_id         (buffer_4_payload_state_id                    ), //i
    .io_inputs_4_payload_state_element    (buffer_4_payload_state_element               ), //i
    .io_inputs_5_valid                    (buffer_5_valid                               ), //i
    .io_inputs_5_ready                    (streamMux_7_io_inputs_5_ready                ), //o
    .io_inputs_5_payload_state_id         (buffer_5_payload_state_id                    ), //i
    .io_inputs_5_payload_state_element    (buffer_5_payload_state_element               ), //i
    .io_output_valid                      (streamMux_7_io_output_valid                  ), //o
    .io_output_ready                      (streamMux_7_io_output_ready                  ), //i
    .io_output_payload_state_id           (streamMux_7_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamMux_7_io_output_payload_state_element  )  //o
  );
  assign when_AXI4StreamInterface_l211 = (io_output_valid && io_output_ready);
  assign _zz_demux_select = {input_demux_5_ready,{input_demux_4_ready,{input_demux_3_ready,{input_demux_2_ready,{input_demux_1_ready,input_demux_0_ready}}}}};
  assign _zz_demux_select_1 = (_zz_demux_select & (~ _zz__zz_demux_select_1));
  assign _zz_demux_select_2 = _zz_demux_select_1[3];
  assign _zz_demux_select_3 = _zz_demux_select_1[5];
  assign _zz_demux_select_4 = ((_zz_demux_select_1[1] || _zz_demux_select_2) || _zz_demux_select_3);
  assign _zz_demux_select_5 = (_zz_demux_select_1[2] || _zz_demux_select_2);
  assign _zz_demux_select_6 = (_zz_demux_select_1[4] || _zz_demux_select_3);
  assign demux_select = {_zz_demux_select_6,{_zz_demux_select_5,_zz_demux_select_4}};
  assign io_input_ready = streamDemux_7_io_input_ready;
  assign input_demux_0_valid = streamDemux_7_io_outputs_0_valid;
  assign input_demux_0_payload_state_id = streamDemux_7_io_outputs_0_payload_state_id;
  assign input_demux_0_payload_state_element = streamDemux_7_io_outputs_0_payload_state_element;
  assign input_demux_1_valid = streamDemux_7_io_outputs_1_valid;
  assign input_demux_1_payload_state_id = streamDemux_7_io_outputs_1_payload_state_id;
  assign input_demux_1_payload_state_element = streamDemux_7_io_outputs_1_payload_state_element;
  assign input_demux_2_valid = streamDemux_7_io_outputs_2_valid;
  assign input_demux_2_payload_state_id = streamDemux_7_io_outputs_2_payload_state_id;
  assign input_demux_2_payload_state_element = streamDemux_7_io_outputs_2_payload_state_element;
  assign input_demux_3_valid = streamDemux_7_io_outputs_3_valid;
  assign input_demux_3_payload_state_id = streamDemux_7_io_outputs_3_payload_state_id;
  assign input_demux_3_payload_state_element = streamDemux_7_io_outputs_3_payload_state_element;
  assign input_demux_4_valid = streamDemux_7_io_outputs_4_valid;
  assign input_demux_4_payload_state_id = streamDemux_7_io_outputs_4_payload_state_id;
  assign input_demux_4_payload_state_element = streamDemux_7_io_outputs_4_payload_state_element;
  assign input_demux_5_valid = streamDemux_7_io_outputs_5_valid;
  assign input_demux_5_payload_state_id = streamDemux_7_io_outputs_5_payload_state_id;
  assign input_demux_5_payload_state_element = streamDemux_7_io_outputs_5_payload_state_element;
  always @(*) begin
    input_demux_0_ready = buffer_0_ready;
    if(when_Stream_l342) begin
      input_demux_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! buffer_0_valid);
  assign buffer_0_valid = input_demux_0_rValid;
  assign buffer_0_payload_state_id = input_demux_0_rData_state_id;
  assign buffer_0_payload_state_element = input_demux_0_rData_state_element;
  always @(*) begin
    input_demux_1_ready = buffer_1_ready;
    if(when_Stream_l342_1) begin
      input_demux_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! buffer_1_valid);
  assign buffer_1_valid = input_demux_1_rValid;
  assign buffer_1_payload_state_id = input_demux_1_rData_state_id;
  assign buffer_1_payload_state_element = input_demux_1_rData_state_element;
  always @(*) begin
    input_demux_2_ready = buffer_2_ready;
    if(when_Stream_l342_2) begin
      input_demux_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! buffer_2_valid);
  assign buffer_2_valid = input_demux_2_rValid;
  assign buffer_2_payload_state_id = input_demux_2_rData_state_id;
  assign buffer_2_payload_state_element = input_demux_2_rData_state_element;
  always @(*) begin
    input_demux_3_ready = buffer_3_ready;
    if(when_Stream_l342_3) begin
      input_demux_3_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! buffer_3_valid);
  assign buffer_3_valid = input_demux_3_rValid;
  assign buffer_3_payload_state_id = input_demux_3_rData_state_id;
  assign buffer_3_payload_state_element = input_demux_3_rData_state_element;
  always @(*) begin
    input_demux_4_ready = buffer_4_ready;
    if(when_Stream_l342_4) begin
      input_demux_4_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! buffer_4_valid);
  assign buffer_4_valid = input_demux_4_rValid;
  assign buffer_4_payload_state_id = input_demux_4_rData_state_id;
  assign buffer_4_payload_state_element = input_demux_4_rData_state_element;
  always @(*) begin
    input_demux_5_ready = buffer_5_ready;
    if(when_Stream_l342_5) begin
      input_demux_5_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! buffer_5_valid);
  assign buffer_5_valid = input_demux_5_rValid;
  assign buffer_5_payload_state_id = input_demux_5_rData_state_id;
  assign buffer_5_payload_state_element = input_demux_5_rData_state_element;
  assign _zz_select = (buffer_3_valid && (buffer_3_payload_state_id == idCounter));
  assign _zz_select_1 = (buffer_5_valid && (buffer_5_payload_state_id == idCounter));
  assign _zz_select_2 = (((buffer_1_valid && (buffer_1_payload_state_id == idCounter)) || _zz_select) || _zz_select_1);
  assign _zz_select_3 = ((buffer_2_valid && (buffer_2_payload_state_id == idCounter)) || _zz_select);
  assign _zz_select_4 = ((buffer_4_valid && (buffer_4_payload_state_id == idCounter)) || _zz_select_1);
  assign select_1 = {_zz_select_4,{_zz_select_3,_zz_select_2}};
  assign buffer_0_ready = streamMux_7_io_inputs_0_ready;
  assign buffer_1_ready = streamMux_7_io_inputs_1_ready;
  assign buffer_2_ready = streamMux_7_io_inputs_2_ready;
  assign buffer_3_ready = streamMux_7_io_inputs_3_ready;
  assign buffer_4_ready = streamMux_7_io_inputs_4_ready;
  assign buffer_5_ready = streamMux_7_io_inputs_5_ready;
  assign io_output_valid = (streamMux_7_io_output_valid && (streamMux_7_io_output_payload_state_id == idCounter));
  assign io_output_last = 1'b1;
  assign io_output_payload = streamMux_7_io_output_payload_state_element;
  assign streamMux_7_io_output_ready = (io_output_ready && (streamMux_7_io_output_payload_state_id == idCounter));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      idCounter <= 7'h0;
      input_demux_0_rValid <= 1'b0;
      input_demux_1_rValid <= 1'b0;
      input_demux_2_rValid <= 1'b0;
      input_demux_3_rValid <= 1'b0;
      input_demux_4_rValid <= 1'b0;
      input_demux_5_rValid <= 1'b0;
    end else begin
      if(when_AXI4StreamInterface_l211) begin
        idCounter <= (idCounter + 7'h01);
      end
      if(input_demux_0_ready) begin
        input_demux_0_rValid <= input_demux_0_valid;
      end
      if(input_demux_1_ready) begin
        input_demux_1_rValid <= input_demux_1_valid;
      end
      if(input_demux_2_ready) begin
        input_demux_2_rValid <= input_demux_2_valid;
      end
      if(input_demux_3_ready) begin
        input_demux_3_rValid <= input_demux_3_valid;
      end
      if(input_demux_4_ready) begin
        input_demux_4_rValid <= input_demux_4_valid;
      end
      if(input_demux_5_ready) begin
        input_demux_5_rValid <= input_demux_5_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(input_demux_0_ready) begin
      input_demux_0_rData_state_id <= input_demux_0_payload_state_id;
      input_demux_0_rData_state_element <= input_demux_0_payload_state_element;
    end
    if(input_demux_1_ready) begin
      input_demux_1_rData_state_id <= input_demux_1_payload_state_id;
      input_demux_1_rData_state_element <= input_demux_1_payload_state_element;
    end
    if(input_demux_2_ready) begin
      input_demux_2_rData_state_id <= input_demux_2_payload_state_id;
      input_demux_2_rData_state_element <= input_demux_2_payload_state_element;
    end
    if(input_demux_3_ready) begin
      input_demux_3_rData_state_id <= input_demux_3_payload_state_id;
      input_demux_3_rData_state_element <= input_demux_3_payload_state_element;
    end
    if(input_demux_4_ready) begin
      input_demux_4_rData_state_id <= input_demux_4_payload_state_id;
      input_demux_4_rData_state_element <= input_demux_4_payload_state_element;
    end
    if(input_demux_5_ready) begin
      input_demux_5_rData_state_id <= input_demux_5_payload_state_id;
      input_demux_5_rData_state_element <= input_demux_5_payload_state_element;
    end
  end


endmodule

module DataLoopbackBuffer (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_elements_0,
  input      [254:0]  io_input_payload_state_elements_1,
  input      [254:0]  io_input_payload_state_elements_2,
  input      [254:0]  io_input_payload_state_elements_3,
  input      [254:0]  io_input_payload_state_elements_4,
  input      [254:0]  io_input_payload_state_elements_5,
  input      [254:0]  io_input_payload_state_elements_6,
  input      [254:0]  io_input_payload_state_elements_7,
  input      [254:0]  io_input_payload_state_elements_8,
  input      [254:0]  io_input_payload_state_elements_9,
  input      [254:0]  io_input_payload_state_elements_10,
  input      [254:0]  io_input_payload_state_elements_11,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_round_index,
  output     [3:0]    io_outputs_0_payload_state_index,
  output     [3:0]    io_outputs_0_payload_state_size,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [254:0]  io_outputs_0_payload_state_element,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_round_index,
  output     [3:0]    io_outputs_1_payload_state_index,
  output     [3:0]    io_outputs_1_payload_state_size,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [254:0]  io_outputs_1_payload_state_element,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [6:0]    io_outputs_2_payload_round_index,
  output     [3:0]    io_outputs_2_payload_state_index,
  output     [3:0]    io_outputs_2_payload_state_size,
  output     [6:0]    io_outputs_2_payload_state_id,
  output     [254:0]  io_outputs_2_payload_state_element,
  output reg [3:0]    io_residue,
  input               clk,
  input               reset
);
  reg                 streamArbiter_12_io_output_ready;
  reg                 streamArbiter_13_io_output_ready;
  reg                 streamArbiter_14_io_output_ready;
  reg                 streamArbiter_15_io_output_ready;
  reg                 streamArbiter_16_io_output_ready;
  reg                 streamArbiter_17_io_output_ready;
  reg                 streamArbiter_18_io_output_ready;
  reg                 streamArbiter_19_io_output_ready;
  reg                 streamArbiter_20_io_output_ready;
  wire                streamArbiter_12_io_inputs_0_ready;
  wire                streamArbiter_12_io_inputs_1_ready;
  wire                streamArbiter_12_io_output_valid;
  wire       [6:0]    streamArbiter_12_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_12_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_12_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_12_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_12_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_12_io_chosen;
  wire       [1:0]    streamArbiter_12_io_chosenOH;
  wire                streamArbiter_13_io_inputs_0_ready;
  wire                streamArbiter_13_io_inputs_1_ready;
  wire                streamArbiter_13_io_output_valid;
  wire       [6:0]    streamArbiter_13_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_13_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_13_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_13_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_13_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_13_io_chosen;
  wire       [1:0]    streamArbiter_13_io_chosenOH;
  wire                streamArbiter_14_io_inputs_0_ready;
  wire                streamArbiter_14_io_inputs_1_ready;
  wire                streamArbiter_14_io_output_valid;
  wire       [6:0]    streamArbiter_14_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_14_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_14_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_14_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_14_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_14_io_chosen;
  wire       [1:0]    streamArbiter_14_io_chosenOH;
  wire                streamArbiter_15_io_inputs_0_ready;
  wire                streamArbiter_15_io_inputs_1_ready;
  wire                streamArbiter_15_io_output_valid;
  wire       [6:0]    streamArbiter_15_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_15_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_15_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_15_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_15_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_15_io_chosen;
  wire       [1:0]    streamArbiter_15_io_chosenOH;
  wire                streamArbiter_16_io_inputs_0_ready;
  wire                streamArbiter_16_io_inputs_1_ready;
  wire                streamArbiter_16_io_output_valid;
  wire       [6:0]    streamArbiter_16_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_16_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_16_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_16_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_16_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_16_io_chosen;
  wire       [1:0]    streamArbiter_16_io_chosenOH;
  wire                streamArbiter_17_io_inputs_0_ready;
  wire                streamArbiter_17_io_inputs_1_ready;
  wire                streamArbiter_17_io_output_valid;
  wire       [6:0]    streamArbiter_17_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_17_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_17_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_17_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_17_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_17_io_chosen;
  wire       [1:0]    streamArbiter_17_io_chosenOH;
  wire                streamArbiter_18_io_inputs_0_ready;
  wire                streamArbiter_18_io_inputs_1_ready;
  wire                streamArbiter_18_io_output_valid;
  wire       [6:0]    streamArbiter_18_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_18_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_18_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_18_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_18_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_18_io_chosen;
  wire       [1:0]    streamArbiter_18_io_chosenOH;
  wire                streamArbiter_19_io_inputs_0_ready;
  wire                streamArbiter_19_io_inputs_1_ready;
  wire                streamArbiter_19_io_output_valid;
  wire       [6:0]    streamArbiter_19_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_19_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_19_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_19_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_19_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_19_io_chosen;
  wire       [1:0]    streamArbiter_19_io_chosenOH;
  wire                streamArbiter_20_io_inputs_0_ready;
  wire                streamArbiter_20_io_inputs_1_ready;
  wire                streamArbiter_20_io_output_valid;
  wire       [6:0]    streamArbiter_20_io_output_payload_round_index;
  wire       [3:0]    streamArbiter_20_io_output_payload_state_index;
  wire       [3:0]    streamArbiter_20_io_output_payload_state_size;
  wire       [6:0]    streamArbiter_20_io_output_payload_state_id;
  wire       [254:0]  streamArbiter_20_io_output_payload_state_element;
  wire       [0:0]    streamArbiter_20_io_chosen;
  wire       [1:0]    streamArbiter_20_io_chosenOH;
  wire       [0:0]    _zz_io_input_ready;
  wire       [1:0]    _zz_io_input_ready_1;
  wire                buffer0_0_valid;
  wire                buffer0_0_ready;
  wire       [6:0]    buffer0_0_payload_round_index;
  wire       [3:0]    buffer0_0_payload_state_index;
  wire       [3:0]    buffer0_0_payload_state_size;
  wire       [6:0]    buffer0_0_payload_state_id;
  wire       [254:0]  buffer0_0_payload_state_element;
  wire                buffer0_1_valid;
  wire                buffer0_1_ready;
  wire       [6:0]    buffer0_1_payload_round_index;
  wire       [3:0]    buffer0_1_payload_state_index;
  wire       [3:0]    buffer0_1_payload_state_size;
  wire       [6:0]    buffer0_1_payload_state_id;
  wire       [254:0]  buffer0_1_payload_state_element;
  wire                buffer0_2_valid;
  wire                buffer0_2_ready;
  wire       [6:0]    buffer0_2_payload_round_index;
  wire       [3:0]    buffer0_2_payload_state_index;
  wire       [3:0]    buffer0_2_payload_state_size;
  wire       [6:0]    buffer0_2_payload_state_id;
  wire       [254:0]  buffer0_2_payload_state_element;
  wire                buffer1_0_valid;
  wire                buffer1_0_ready;
  wire       [6:0]    buffer1_0_payload_round_index;
  wire       [3:0]    buffer1_0_payload_state_index;
  wire       [3:0]    buffer1_0_payload_state_size;
  wire       [6:0]    buffer1_0_payload_state_id;
  wire       [254:0]  buffer1_0_payload_state_element;
  wire                buffer1_1_valid;
  wire                buffer1_1_ready;
  wire       [6:0]    buffer1_1_payload_round_index;
  wire       [3:0]    buffer1_1_payload_state_index;
  wire       [3:0]    buffer1_1_payload_state_size;
  wire       [6:0]    buffer1_1_payload_state_id;
  wire       [254:0]  buffer1_1_payload_state_element;
  wire                buffer1_2_valid;
  wire                buffer1_2_ready;
  wire       [6:0]    buffer1_2_payload_round_index;
  wire       [3:0]    buffer1_2_payload_state_index;
  wire       [3:0]    buffer1_2_payload_state_size;
  wire       [6:0]    buffer1_2_payload_state_id;
  wire       [254:0]  buffer1_2_payload_state_element;
  wire                buffer2_0_valid;
  wire                buffer2_0_ready;
  wire       [6:0]    buffer2_0_payload_round_index;
  wire       [3:0]    buffer2_0_payload_state_index;
  wire       [3:0]    buffer2_0_payload_state_size;
  wire       [6:0]    buffer2_0_payload_state_id;
  wire       [254:0]  buffer2_0_payload_state_element;
  wire                buffer2_1_valid;
  wire                buffer2_1_ready;
  wire       [6:0]    buffer2_1_payload_round_index;
  wire       [3:0]    buffer2_1_payload_state_index;
  wire       [3:0]    buffer2_1_payload_state_size;
  wire       [6:0]    buffer2_1_payload_state_id;
  wire       [254:0]  buffer2_1_payload_state_element;
  wire                buffer2_2_valid;
  wire                buffer2_2_ready;
  wire       [6:0]    buffer2_2_payload_round_index;
  wire       [3:0]    buffer2_2_payload_state_index;
  wire       [3:0]    buffer2_2_payload_state_size;
  wire       [6:0]    buffer2_2_payload_state_id;
  wire       [254:0]  buffer2_2_payload_state_element;
  wire                buffer3_0_valid;
  reg                 buffer3_0_ready;
  wire       [6:0]    buffer3_0_payload_round_index;
  wire       [3:0]    buffer3_0_payload_state_index;
  wire       [3:0]    buffer3_0_payload_state_size;
  wire       [6:0]    buffer3_0_payload_state_id;
  wire       [254:0]  buffer3_0_payload_state_element;
  wire                buffer3_1_valid;
  reg                 buffer3_1_ready;
  wire       [6:0]    buffer3_1_payload_round_index;
  wire       [3:0]    buffer3_1_payload_state_index;
  wire       [3:0]    buffer3_1_payload_state_size;
  wire       [6:0]    buffer3_1_payload_state_id;
  wire       [254:0]  buffer3_1_payload_state_element;
  wire                buffer3_2_valid;
  reg                 buffer3_2_ready;
  wire       [6:0]    buffer3_2_payload_round_index;
  wire       [3:0]    buffer3_2_payload_state_index;
  wire       [3:0]    buffer3_2_payload_state_size;
  wire       [6:0]    buffer3_2_payload_state_id;
  wire       [254:0]  buffer3_2_payload_state_element;
  wire                inputs_0_valid;
  reg                 inputs_0_ready;
  wire       [6:0]    inputs_0_payload_round_index;
  wire       [3:0]    inputs_0_payload_state_index;
  wire       [3:0]    inputs_0_payload_state_size;
  wire       [6:0]    inputs_0_payload_state_id;
  wire       [254:0]  inputs_0_payload_state_element;
  wire                inputs_1_valid;
  reg                 inputs_1_ready;
  wire       [6:0]    inputs_1_payload_round_index;
  wire       [3:0]    inputs_1_payload_state_index;
  wire       [3:0]    inputs_1_payload_state_size;
  wire       [6:0]    inputs_1_payload_state_id;
  wire       [254:0]  inputs_1_payload_state_element;
  wire                inputs_2_valid;
  reg                 inputs_2_ready;
  wire       [6:0]    inputs_2_payload_round_index;
  wire       [3:0]    inputs_2_payload_state_index;
  wire       [3:0]    inputs_2_payload_state_size;
  wire       [6:0]    inputs_2_payload_state_id;
  wire       [254:0]  inputs_2_payload_state_element;
  wire                inputs_3_valid;
  reg                 inputs_3_ready;
  wire       [6:0]    inputs_3_payload_round_index;
  wire       [3:0]    inputs_3_payload_state_index;
  wire       [3:0]    inputs_3_payload_state_size;
  wire       [6:0]    inputs_3_payload_state_id;
  wire       [254:0]  inputs_3_payload_state_element;
  wire                inputs_4_valid;
  reg                 inputs_4_ready;
  wire       [6:0]    inputs_4_payload_round_index;
  wire       [3:0]    inputs_4_payload_state_index;
  wire       [3:0]    inputs_4_payload_state_size;
  wire       [6:0]    inputs_4_payload_state_id;
  wire       [254:0]  inputs_4_payload_state_element;
  wire                inputs_5_valid;
  reg                 inputs_5_ready;
  wire       [6:0]    inputs_5_payload_round_index;
  wire       [3:0]    inputs_5_payload_state_index;
  wire       [3:0]    inputs_5_payload_state_size;
  wire       [6:0]    inputs_5_payload_state_id;
  wire       [254:0]  inputs_5_payload_state_element;
  wire                inputs_6_valid;
  reg                 inputs_6_ready;
  wire       [6:0]    inputs_6_payload_round_index;
  wire       [3:0]    inputs_6_payload_state_index;
  wire       [3:0]    inputs_6_payload_state_size;
  wire       [6:0]    inputs_6_payload_state_id;
  wire       [254:0]  inputs_6_payload_state_element;
  wire                inputs_7_valid;
  reg                 inputs_7_ready;
  wire       [6:0]    inputs_7_payload_round_index;
  wire       [3:0]    inputs_7_payload_state_index;
  wire       [3:0]    inputs_7_payload_state_size;
  wire       [6:0]    inputs_7_payload_state_id;
  wire       [254:0]  inputs_7_payload_state_element;
  wire                inputs_8_valid;
  reg                 inputs_8_ready;
  wire       [6:0]    inputs_8_payload_round_index;
  wire       [3:0]    inputs_8_payload_state_index;
  wire       [3:0]    inputs_8_payload_state_size;
  wire       [6:0]    inputs_8_payload_state_id;
  wire       [254:0]  inputs_8_payload_state_element;
  wire                inputs_9_valid;
  reg                 inputs_9_ready;
  wire       [6:0]    inputs_9_payload_round_index;
  wire       [3:0]    inputs_9_payload_state_index;
  wire       [3:0]    inputs_9_payload_state_size;
  wire       [6:0]    inputs_9_payload_state_id;
  wire       [254:0]  inputs_9_payload_state_element;
  wire                inputs_10_valid;
  reg                 inputs_10_ready;
  wire       [6:0]    inputs_10_payload_round_index;
  wire       [3:0]    inputs_10_payload_state_index;
  wire       [3:0]    inputs_10_payload_state_size;
  wire       [6:0]    inputs_10_payload_state_id;
  wire       [254:0]  inputs_10_payload_state_element;
  wire                inputs_11_valid;
  reg                 inputs_11_ready;
  wire       [6:0]    inputs_11_payload_round_index;
  wire       [3:0]    inputs_11_payload_state_index;
  wire       [3:0]    inputs_11_payload_state_size;
  wire       [6:0]    inputs_11_payload_state_id;
  wire       [254:0]  inputs_11_payload_state_element;
  wire                inputs_0_m2sPipe_valid;
  wire                inputs_0_m2sPipe_ready;
  wire       [6:0]    inputs_0_m2sPipe_payload_round_index;
  wire       [3:0]    inputs_0_m2sPipe_payload_state_index;
  wire       [3:0]    inputs_0_m2sPipe_payload_state_size;
  wire       [6:0]    inputs_0_m2sPipe_payload_state_id;
  wire       [254:0]  inputs_0_m2sPipe_payload_state_element;
  reg                 inputs_0_rValid;
  reg        [6:0]    inputs_0_rData_round_index;
  reg        [3:0]    inputs_0_rData_state_index;
  reg        [3:0]    inputs_0_rData_state_size;
  reg        [6:0]    inputs_0_rData_state_id;
  reg        [254:0]  inputs_0_rData_state_element;
  wire                when_Stream_l342;
  wire                when_Stream_l408;
  reg                 inputs_3_thrown_valid;
  wire                inputs_3_thrown_ready;
  wire       [6:0]    inputs_3_thrown_payload_round_index;
  wire       [3:0]    inputs_3_thrown_payload_state_index;
  wire       [3:0]    inputs_3_thrown_payload_state_size;
  wire       [6:0]    inputs_3_thrown_payload_state_id;
  wire       [254:0]  inputs_3_thrown_payload_state_element;
  wire                streamArbiter_12_io_output_m2sPipe_valid;
  wire                streamArbiter_12_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_12_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_12_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_12_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_12_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_12_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_12_io_output_rValid;
  reg        [6:0]    streamArbiter_12_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_12_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_12_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_12_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_12_io_output_rData_state_element;
  wire                when_Stream_l342_1;
  wire                when_Stream_l408_1;
  reg                 inputs_6_thrown_valid;
  wire                inputs_6_thrown_ready;
  wire       [6:0]    inputs_6_thrown_payload_round_index;
  wire       [3:0]    inputs_6_thrown_payload_state_index;
  wire       [3:0]    inputs_6_thrown_payload_state_size;
  wire       [6:0]    inputs_6_thrown_payload_state_id;
  wire       [254:0]  inputs_6_thrown_payload_state_element;
  wire                streamArbiter_13_io_output_m2sPipe_valid;
  wire                streamArbiter_13_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_13_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_13_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_13_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_13_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_13_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_13_io_output_rValid;
  reg        [6:0]    streamArbiter_13_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_13_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_13_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_13_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_13_io_output_rData_state_element;
  wire                when_Stream_l342_2;
  wire                when_Stream_l408_2;
  reg                 inputs_9_thrown_valid;
  wire                inputs_9_thrown_ready;
  wire       [6:0]    inputs_9_thrown_payload_round_index;
  wire       [3:0]    inputs_9_thrown_payload_state_index;
  wire       [3:0]    inputs_9_thrown_payload_state_size;
  wire       [6:0]    inputs_9_thrown_payload_state_id;
  wire       [254:0]  inputs_9_thrown_payload_state_element;
  wire                streamArbiter_14_io_output_m2sPipe_valid;
  wire                streamArbiter_14_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_14_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_14_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_14_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_14_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_14_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_14_io_output_rValid;
  reg        [6:0]    streamArbiter_14_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_14_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_14_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_14_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_14_io_output_rData_state_element;
  wire                when_Stream_l342_3;
  wire                inputs_1_m2sPipe_valid;
  wire                inputs_1_m2sPipe_ready;
  wire       [6:0]    inputs_1_m2sPipe_payload_round_index;
  wire       [3:0]    inputs_1_m2sPipe_payload_state_index;
  wire       [3:0]    inputs_1_m2sPipe_payload_state_size;
  wire       [6:0]    inputs_1_m2sPipe_payload_state_id;
  wire       [254:0]  inputs_1_m2sPipe_payload_state_element;
  reg                 inputs_1_rValid;
  reg        [6:0]    inputs_1_rData_round_index;
  reg        [3:0]    inputs_1_rData_state_index;
  reg        [3:0]    inputs_1_rData_state_size;
  reg        [6:0]    inputs_1_rData_state_id;
  reg        [254:0]  inputs_1_rData_state_element;
  wire                when_Stream_l342_4;
  wire                when_Stream_l408_3;
  reg                 inputs_4_thrown_valid;
  wire                inputs_4_thrown_ready;
  wire       [6:0]    inputs_4_thrown_payload_round_index;
  wire       [3:0]    inputs_4_thrown_payload_state_index;
  wire       [3:0]    inputs_4_thrown_payload_state_size;
  wire       [6:0]    inputs_4_thrown_payload_state_id;
  wire       [254:0]  inputs_4_thrown_payload_state_element;
  wire                streamArbiter_15_io_output_m2sPipe_valid;
  wire                streamArbiter_15_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_15_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_15_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_15_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_15_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_15_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_15_io_output_rValid;
  reg        [6:0]    streamArbiter_15_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_15_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_15_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_15_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_15_io_output_rData_state_element;
  wire                when_Stream_l342_5;
  wire                when_Stream_l408_4;
  reg                 inputs_7_thrown_valid;
  wire                inputs_7_thrown_ready;
  wire       [6:0]    inputs_7_thrown_payload_round_index;
  wire       [3:0]    inputs_7_thrown_payload_state_index;
  wire       [3:0]    inputs_7_thrown_payload_state_size;
  wire       [6:0]    inputs_7_thrown_payload_state_id;
  wire       [254:0]  inputs_7_thrown_payload_state_element;
  wire                streamArbiter_16_io_output_m2sPipe_valid;
  wire                streamArbiter_16_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_16_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_16_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_16_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_16_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_16_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_16_io_output_rValid;
  reg        [6:0]    streamArbiter_16_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_16_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_16_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_16_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_16_io_output_rData_state_element;
  wire                when_Stream_l342_6;
  wire                when_Stream_l408_5;
  reg                 inputs_10_thrown_valid;
  wire                inputs_10_thrown_ready;
  wire       [6:0]    inputs_10_thrown_payload_round_index;
  wire       [3:0]    inputs_10_thrown_payload_state_index;
  wire       [3:0]    inputs_10_thrown_payload_state_size;
  wire       [6:0]    inputs_10_thrown_payload_state_id;
  wire       [254:0]  inputs_10_thrown_payload_state_element;
  wire                streamArbiter_17_io_output_m2sPipe_valid;
  wire                streamArbiter_17_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_17_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_17_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_17_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_17_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_17_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_17_io_output_rValid;
  reg        [6:0]    streamArbiter_17_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_17_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_17_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_17_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_17_io_output_rData_state_element;
  wire                when_Stream_l342_7;
  wire                inputs_2_m2sPipe_valid;
  wire                inputs_2_m2sPipe_ready;
  wire       [6:0]    inputs_2_m2sPipe_payload_round_index;
  wire       [3:0]    inputs_2_m2sPipe_payload_state_index;
  wire       [3:0]    inputs_2_m2sPipe_payload_state_size;
  wire       [6:0]    inputs_2_m2sPipe_payload_state_id;
  wire       [254:0]  inputs_2_m2sPipe_payload_state_element;
  reg                 inputs_2_rValid;
  reg        [6:0]    inputs_2_rData_round_index;
  reg        [3:0]    inputs_2_rData_state_index;
  reg        [3:0]    inputs_2_rData_state_size;
  reg        [6:0]    inputs_2_rData_state_id;
  reg        [254:0]  inputs_2_rData_state_element;
  wire                when_Stream_l342_8;
  wire                when_Stream_l408_6;
  reg                 inputs_5_thrown_valid;
  wire                inputs_5_thrown_ready;
  wire       [6:0]    inputs_5_thrown_payload_round_index;
  wire       [3:0]    inputs_5_thrown_payload_state_index;
  wire       [3:0]    inputs_5_thrown_payload_state_size;
  wire       [6:0]    inputs_5_thrown_payload_state_id;
  wire       [254:0]  inputs_5_thrown_payload_state_element;
  wire                streamArbiter_18_io_output_m2sPipe_valid;
  wire                streamArbiter_18_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_18_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_18_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_18_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_18_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_18_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_18_io_output_rValid;
  reg        [6:0]    streamArbiter_18_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_18_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_18_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_18_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_18_io_output_rData_state_element;
  wire                when_Stream_l342_9;
  wire                when_Stream_l408_7;
  reg                 inputs_8_thrown_valid;
  wire                inputs_8_thrown_ready;
  wire       [6:0]    inputs_8_thrown_payload_round_index;
  wire       [3:0]    inputs_8_thrown_payload_state_index;
  wire       [3:0]    inputs_8_thrown_payload_state_size;
  wire       [6:0]    inputs_8_thrown_payload_state_id;
  wire       [254:0]  inputs_8_thrown_payload_state_element;
  wire                streamArbiter_19_io_output_m2sPipe_valid;
  wire                streamArbiter_19_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_19_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_19_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_19_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_19_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_19_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_19_io_output_rValid;
  reg        [6:0]    streamArbiter_19_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_19_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_19_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_19_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_19_io_output_rData_state_element;
  wire                when_Stream_l342_10;
  wire                when_Stream_l408_8;
  reg                 inputs_11_thrown_valid;
  wire                inputs_11_thrown_ready;
  wire       [6:0]    inputs_11_thrown_payload_round_index;
  wire       [3:0]    inputs_11_thrown_payload_state_index;
  wire       [3:0]    inputs_11_thrown_payload_state_size;
  wire       [6:0]    inputs_11_thrown_payload_state_id;
  wire       [254:0]  inputs_11_thrown_payload_state_element;
  wire                streamArbiter_20_io_output_m2sPipe_valid;
  wire                streamArbiter_20_io_output_m2sPipe_ready;
  wire       [6:0]    streamArbiter_20_io_output_m2sPipe_payload_round_index;
  wire       [3:0]    streamArbiter_20_io_output_m2sPipe_payload_state_index;
  wire       [3:0]    streamArbiter_20_io_output_m2sPipe_payload_state_size;
  wire       [6:0]    streamArbiter_20_io_output_m2sPipe_payload_state_id;
  wire       [254:0]  streamArbiter_20_io_output_m2sPipe_payload_state_element;
  reg                 streamArbiter_20_io_output_rValid;
  reg        [6:0]    streamArbiter_20_io_output_rData_round_index;
  reg        [3:0]    streamArbiter_20_io_output_rData_state_index;
  reg        [3:0]    streamArbiter_20_io_output_rData_state_size;
  reg        [6:0]    streamArbiter_20_io_output_rData_state_id;
  reg        [254:0]  streamArbiter_20_io_output_rData_state_element;
  wire                when_Stream_l342_11;
  wire                buffers_0_0_valid;
  reg                 buffers_0_0_ready;
  wire       [6:0]    buffers_0_0_payload_round_index;
  wire       [3:0]    buffers_0_0_payload_state_index;
  wire       [3:0]    buffers_0_0_payload_state_size;
  wire       [6:0]    buffers_0_0_payload_state_id;
  wire       [254:0]  buffers_0_0_payload_state_element;
  wire                buffers_0_1_valid;
  reg                 buffers_0_1_ready;
  wire       [6:0]    buffers_0_1_payload_round_index;
  wire       [3:0]    buffers_0_1_payload_state_index;
  wire       [3:0]    buffers_0_1_payload_state_size;
  wire       [6:0]    buffers_0_1_payload_state_id;
  wire       [254:0]  buffers_0_1_payload_state_element;
  wire                buffers_0_2_valid;
  reg                 buffers_0_2_ready;
  wire       [6:0]    buffers_0_2_payload_round_index;
  wire       [3:0]    buffers_0_2_payload_state_index;
  wire       [3:0]    buffers_0_2_payload_state_size;
  wire       [6:0]    buffers_0_2_payload_state_id;
  wire       [254:0]  buffers_0_2_payload_state_element;
  wire                buffers_1_0_valid;
  reg                 buffers_1_0_ready;
  wire       [6:0]    buffers_1_0_payload_round_index;
  wire       [3:0]    buffers_1_0_payload_state_index;
  wire       [3:0]    buffers_1_0_payload_state_size;
  wire       [6:0]    buffers_1_0_payload_state_id;
  wire       [254:0]  buffers_1_0_payload_state_element;
  wire                buffers_1_1_valid;
  reg                 buffers_1_1_ready;
  wire       [6:0]    buffers_1_1_payload_round_index;
  wire       [3:0]    buffers_1_1_payload_state_index;
  wire       [3:0]    buffers_1_1_payload_state_size;
  wire       [6:0]    buffers_1_1_payload_state_id;
  wire       [254:0]  buffers_1_1_payload_state_element;
  wire                buffers_1_2_valid;
  reg                 buffers_1_2_ready;
  wire       [6:0]    buffers_1_2_payload_round_index;
  wire       [3:0]    buffers_1_2_payload_state_index;
  wire       [3:0]    buffers_1_2_payload_state_size;
  wire       [6:0]    buffers_1_2_payload_state_id;
  wire       [254:0]  buffers_1_2_payload_state_element;
  wire                buffers_2_0_valid;
  reg                 buffers_2_0_ready;
  wire       [6:0]    buffers_2_0_payload_round_index;
  wire       [3:0]    buffers_2_0_payload_state_index;
  wire       [3:0]    buffers_2_0_payload_state_size;
  wire       [6:0]    buffers_2_0_payload_state_id;
  wire       [254:0]  buffers_2_0_payload_state_element;
  wire                buffers_2_1_valid;
  reg                 buffers_2_1_ready;
  wire       [6:0]    buffers_2_1_payload_round_index;
  wire       [3:0]    buffers_2_1_payload_state_index;
  wire       [3:0]    buffers_2_1_payload_state_size;
  wire       [6:0]    buffers_2_1_payload_state_id;
  wire       [254:0]  buffers_2_1_payload_state_element;
  wire                buffers_2_2_valid;
  reg                 buffers_2_2_ready;
  wire       [6:0]    buffers_2_2_payload_round_index;
  wire       [3:0]    buffers_2_2_payload_state_index;
  wire       [3:0]    buffers_2_2_payload_state_size;
  wire       [6:0]    buffers_2_2_payload_state_id;
  wire       [254:0]  buffers_2_2_payload_state_element;
  wire                buffers_3_0_valid;
  wire                buffers_3_0_ready;
  wire       [6:0]    buffers_3_0_payload_round_index;
  wire       [3:0]    buffers_3_0_payload_state_index;
  wire       [3:0]    buffers_3_0_payload_state_size;
  wire       [6:0]    buffers_3_0_payload_state_id;
  wire       [254:0]  buffers_3_0_payload_state_element;
  wire                buffers_3_1_valid;
  wire                buffers_3_1_ready;
  wire       [6:0]    buffers_3_1_payload_round_index;
  wire       [3:0]    buffers_3_1_payload_state_index;
  wire       [3:0]    buffers_3_1_payload_state_size;
  wire       [6:0]    buffers_3_1_payload_state_id;
  wire       [254:0]  buffers_3_1_payload_state_element;
  wire                buffers_3_2_valid;
  wire                buffers_3_2_ready;
  wire       [6:0]    buffers_3_2_payload_round_index;
  wire       [3:0]    buffers_3_2_payload_state_index;
  wire       [3:0]    buffers_3_2_payload_state_size;
  wire       [6:0]    buffers_3_2_payload_state_id;
  wire       [254:0]  buffers_3_2_payload_state_element;
  wire                buffer3_0_m2sPipe_valid;
  wire                buffer3_0_m2sPipe_ready;
  wire       [6:0]    buffer3_0_m2sPipe_payload_round_index;
  wire       [3:0]    buffer3_0_m2sPipe_payload_state_index;
  wire       [3:0]    buffer3_0_m2sPipe_payload_state_size;
  wire       [6:0]    buffer3_0_m2sPipe_payload_state_id;
  wire       [254:0]  buffer3_0_m2sPipe_payload_state_element;
  reg                 buffer3_0_rValid;
  reg        [6:0]    buffer3_0_rData_round_index;
  reg        [3:0]    buffer3_0_rData_state_index;
  reg        [3:0]    buffer3_0_rData_state_size;
  reg        [6:0]    buffer3_0_rData_state_id;
  reg        [254:0]  buffer3_0_rData_state_element;
  wire                when_Stream_l342_12;
  wire                buffer3_1_m2sPipe_valid;
  wire                buffer3_1_m2sPipe_ready;
  wire       [6:0]    buffer3_1_m2sPipe_payload_round_index;
  wire       [3:0]    buffer3_1_m2sPipe_payload_state_index;
  wire       [3:0]    buffer3_1_m2sPipe_payload_state_size;
  wire       [6:0]    buffer3_1_m2sPipe_payload_state_id;
  wire       [254:0]  buffer3_1_m2sPipe_payload_state_element;
  reg                 buffer3_1_rValid;
  reg        [6:0]    buffer3_1_rData_round_index;
  reg        [3:0]    buffer3_1_rData_state_index;
  reg        [3:0]    buffer3_1_rData_state_size;
  reg        [6:0]    buffer3_1_rData_state_id;
  reg        [254:0]  buffer3_1_rData_state_element;
  wire                when_Stream_l342_13;
  wire                buffer3_2_m2sPipe_valid;
  wire                buffer3_2_m2sPipe_ready;
  wire       [6:0]    buffer3_2_m2sPipe_payload_round_index;
  wire       [3:0]    buffer3_2_m2sPipe_payload_state_index;
  wire       [3:0]    buffer3_2_m2sPipe_payload_state_size;
  wire       [6:0]    buffer3_2_m2sPipe_payload_state_id;
  wire       [254:0]  buffer3_2_m2sPipe_payload_state_element;
  reg                 buffer3_2_rValid;
  reg        [6:0]    buffer3_2_rData_round_index;
  reg        [3:0]    buffer3_2_rData_state_index;
  reg        [3:0]    buffer3_2_rData_state_size;
  reg        [6:0]    buffer3_2_rData_state_id;
  reg        [254:0]  buffer3_2_rData_state_element;
  wire                when_Stream_l342_14;
  wire                buffers_0_0_m2sPipe_valid;
  wire                buffers_0_0_m2sPipe_ready;
  wire       [6:0]    buffers_0_0_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_0_0_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_0_0_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_0_0_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_0_0_m2sPipe_payload_state_element;
  reg                 buffers_0_0_rValid;
  reg        [6:0]    buffers_0_0_rData_round_index;
  reg        [3:0]    buffers_0_0_rData_state_index;
  reg        [3:0]    buffers_0_0_rData_state_size;
  reg        [6:0]    buffers_0_0_rData_state_id;
  reg        [254:0]  buffers_0_0_rData_state_element;
  wire                when_Stream_l342_15;
  wire                buffers_0_1_m2sPipe_valid;
  wire                buffers_0_1_m2sPipe_ready;
  wire       [6:0]    buffers_0_1_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_0_1_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_0_1_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_0_1_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_0_1_m2sPipe_payload_state_element;
  reg                 buffers_0_1_rValid;
  reg        [6:0]    buffers_0_1_rData_round_index;
  reg        [3:0]    buffers_0_1_rData_state_index;
  reg        [3:0]    buffers_0_1_rData_state_size;
  reg        [6:0]    buffers_0_1_rData_state_id;
  reg        [254:0]  buffers_0_1_rData_state_element;
  wire                when_Stream_l342_16;
  wire                buffers_0_2_m2sPipe_valid;
  wire                buffers_0_2_m2sPipe_ready;
  wire       [6:0]    buffers_0_2_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_0_2_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_0_2_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_0_2_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_0_2_m2sPipe_payload_state_element;
  reg                 buffers_0_2_rValid;
  reg        [6:0]    buffers_0_2_rData_round_index;
  reg        [3:0]    buffers_0_2_rData_state_index;
  reg        [3:0]    buffers_0_2_rData_state_size;
  reg        [6:0]    buffers_0_2_rData_state_id;
  reg        [254:0]  buffers_0_2_rData_state_element;
  wire                when_Stream_l342_17;
  wire                buffers_1_0_m2sPipe_valid;
  wire                buffers_1_0_m2sPipe_ready;
  wire       [6:0]    buffers_1_0_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_1_0_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_1_0_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_1_0_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_1_0_m2sPipe_payload_state_element;
  reg                 buffers_1_0_rValid;
  reg        [6:0]    buffers_1_0_rData_round_index;
  reg        [3:0]    buffers_1_0_rData_state_index;
  reg        [3:0]    buffers_1_0_rData_state_size;
  reg        [6:0]    buffers_1_0_rData_state_id;
  reg        [254:0]  buffers_1_0_rData_state_element;
  wire                when_Stream_l342_18;
  wire                buffers_1_1_m2sPipe_valid;
  wire                buffers_1_1_m2sPipe_ready;
  wire       [6:0]    buffers_1_1_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_1_1_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_1_1_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_1_1_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_1_1_m2sPipe_payload_state_element;
  reg                 buffers_1_1_rValid;
  reg        [6:0]    buffers_1_1_rData_round_index;
  reg        [3:0]    buffers_1_1_rData_state_index;
  reg        [3:0]    buffers_1_1_rData_state_size;
  reg        [6:0]    buffers_1_1_rData_state_id;
  reg        [254:0]  buffers_1_1_rData_state_element;
  wire                when_Stream_l342_19;
  wire                buffers_1_2_m2sPipe_valid;
  wire                buffers_1_2_m2sPipe_ready;
  wire       [6:0]    buffers_1_2_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_1_2_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_1_2_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_1_2_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_1_2_m2sPipe_payload_state_element;
  reg                 buffers_1_2_rValid;
  reg        [6:0]    buffers_1_2_rData_round_index;
  reg        [3:0]    buffers_1_2_rData_state_index;
  reg        [3:0]    buffers_1_2_rData_state_size;
  reg        [6:0]    buffers_1_2_rData_state_id;
  reg        [254:0]  buffers_1_2_rData_state_element;
  wire                when_Stream_l342_20;
  wire                buffers_2_0_m2sPipe_valid;
  wire                buffers_2_0_m2sPipe_ready;
  wire       [6:0]    buffers_2_0_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_2_0_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_2_0_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_2_0_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_2_0_m2sPipe_payload_state_element;
  reg                 buffers_2_0_rValid;
  reg        [6:0]    buffers_2_0_rData_round_index;
  reg        [3:0]    buffers_2_0_rData_state_index;
  reg        [3:0]    buffers_2_0_rData_state_size;
  reg        [6:0]    buffers_2_0_rData_state_id;
  reg        [254:0]  buffers_2_0_rData_state_element;
  wire                when_Stream_l342_21;
  wire                buffers_2_1_m2sPipe_valid;
  wire                buffers_2_1_m2sPipe_ready;
  wire       [6:0]    buffers_2_1_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_2_1_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_2_1_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_2_1_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_2_1_m2sPipe_payload_state_element;
  reg                 buffers_2_1_rValid;
  reg        [6:0]    buffers_2_1_rData_round_index;
  reg        [3:0]    buffers_2_1_rData_state_index;
  reg        [3:0]    buffers_2_1_rData_state_size;
  reg        [6:0]    buffers_2_1_rData_state_id;
  reg        [254:0]  buffers_2_1_rData_state_element;
  wire                when_Stream_l342_22;
  wire                buffers_2_2_m2sPipe_valid;
  wire                buffers_2_2_m2sPipe_ready;
  wire       [6:0]    buffers_2_2_m2sPipe_payload_round_index;
  wire       [3:0]    buffers_2_2_m2sPipe_payload_state_index;
  wire       [3:0]    buffers_2_2_m2sPipe_payload_state_size;
  wire       [6:0]    buffers_2_2_m2sPipe_payload_state_id;
  wire       [254:0]  buffers_2_2_m2sPipe_payload_state_element;
  reg                 buffers_2_2_rValid;
  reg        [6:0]    buffers_2_2_rData_round_index;
  reg        [3:0]    buffers_2_2_rData_state_index;
  reg        [3:0]    buffers_2_2_rData_state_size;
  reg        [6:0]    buffers_2_2_rData_state_id;
  reg        [254:0]  buffers_2_2_rData_state_element;
  wire                when_Stream_l342_23;
  wire                when_PoseidonTopLevel_l90;
  wire                when_PoseidonTopLevel_l93;
  wire                when_PoseidonTopLevel_l96;
  wire                when_PoseidonTopLevel_l99;

  assign _zz_io_input_ready = inputs_2_ready;
  assign _zz_io_input_ready_1 = {inputs_1_ready,inputs_0_ready};
  StreamArbiter streamArbiter_12 (
    .io_inputs_0_valid                    (buffer0_0_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_12_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer0_0_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer0_0_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer0_0_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer0_0_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer0_0_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_3_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_12_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_3_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_3_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_3_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_3_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_3_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_12_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_12_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_12_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_12_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_12_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_12_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_12_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_12_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_12_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_13 (
    .io_inputs_0_valid                    (buffer1_0_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_13_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer1_0_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer1_0_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer1_0_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer1_0_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer1_0_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_6_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_13_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_6_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_6_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_6_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_6_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_6_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_13_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_13_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_13_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_13_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_13_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_13_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_13_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_13_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_13_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_14 (
    .io_inputs_0_valid                    (buffer2_0_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_14_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer2_0_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer2_0_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer2_0_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer2_0_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer2_0_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_9_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_14_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_9_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_9_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_9_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_9_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_9_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_14_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_14_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_14_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_14_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_14_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_14_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_14_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_14_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_14_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_15 (
    .io_inputs_0_valid                    (buffer0_1_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_15_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer0_1_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer0_1_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer0_1_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer0_1_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer0_1_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_4_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_15_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_4_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_4_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_4_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_4_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_4_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_15_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_15_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_15_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_15_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_15_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_15_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_15_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_15_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_15_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_16 (
    .io_inputs_0_valid                    (buffer1_1_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_16_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer1_1_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer1_1_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer1_1_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer1_1_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer1_1_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_7_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_16_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_7_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_7_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_7_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_7_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_7_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_16_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_16_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_16_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_16_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_16_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_16_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_16_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_16_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_16_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_17 (
    .io_inputs_0_valid                    (buffer2_1_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_17_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer2_1_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer2_1_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer2_1_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer2_1_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer2_1_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_10_thrown_valid                            ), //i
    .io_inputs_1_ready                    (streamArbiter_17_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_10_thrown_payload_round_index              ), //i
    .io_inputs_1_payload_state_index      (inputs_10_thrown_payload_state_index              ), //i
    .io_inputs_1_payload_state_size       (inputs_10_thrown_payload_state_size               ), //i
    .io_inputs_1_payload_state_id         (inputs_10_thrown_payload_state_id                 ), //i
    .io_inputs_1_payload_state_element    (inputs_10_thrown_payload_state_element            ), //i
    .io_output_valid                      (streamArbiter_17_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_17_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_17_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_17_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_17_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_17_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_17_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_17_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_17_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_18 (
    .io_inputs_0_valid                    (buffer0_2_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_18_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer0_2_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer0_2_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer0_2_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer0_2_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer0_2_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_5_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_18_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_5_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_5_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_5_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_5_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_5_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_18_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_18_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_18_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_18_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_18_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_18_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_18_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_18_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_18_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_19 (
    .io_inputs_0_valid                    (buffer1_2_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_19_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer1_2_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer1_2_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer1_2_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer1_2_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer1_2_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_8_thrown_valid                             ), //i
    .io_inputs_1_ready                    (streamArbiter_19_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_8_thrown_payload_round_index               ), //i
    .io_inputs_1_payload_state_index      (inputs_8_thrown_payload_state_index               ), //i
    .io_inputs_1_payload_state_size       (inputs_8_thrown_payload_state_size                ), //i
    .io_inputs_1_payload_state_id         (inputs_8_thrown_payload_state_id                  ), //i
    .io_inputs_1_payload_state_element    (inputs_8_thrown_payload_state_element             ), //i
    .io_output_valid                      (streamArbiter_19_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_19_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_19_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_19_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_19_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_19_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_19_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_19_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_19_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  StreamArbiter streamArbiter_20 (
    .io_inputs_0_valid                    (buffer2_2_valid                                   ), //i
    .io_inputs_0_ready                    (streamArbiter_20_io_inputs_0_ready                ), //o
    .io_inputs_0_payload_round_index      (buffer2_2_payload_round_index                     ), //i
    .io_inputs_0_payload_state_index      (buffer2_2_payload_state_index                     ), //i
    .io_inputs_0_payload_state_size       (buffer2_2_payload_state_size                      ), //i
    .io_inputs_0_payload_state_id         (buffer2_2_payload_state_id                        ), //i
    .io_inputs_0_payload_state_element    (buffer2_2_payload_state_element                   ), //i
    .io_inputs_1_valid                    (inputs_11_thrown_valid                            ), //i
    .io_inputs_1_ready                    (streamArbiter_20_io_inputs_1_ready                ), //o
    .io_inputs_1_payload_round_index      (inputs_11_thrown_payload_round_index              ), //i
    .io_inputs_1_payload_state_index      (inputs_11_thrown_payload_state_index              ), //i
    .io_inputs_1_payload_state_size       (inputs_11_thrown_payload_state_size               ), //i
    .io_inputs_1_payload_state_id         (inputs_11_thrown_payload_state_id                 ), //i
    .io_inputs_1_payload_state_element    (inputs_11_thrown_payload_state_element            ), //i
    .io_output_valid                      (streamArbiter_20_io_output_valid                  ), //o
    .io_output_ready                      (streamArbiter_20_io_output_ready                  ), //i
    .io_output_payload_round_index        (streamArbiter_20_io_output_payload_round_index    ), //o
    .io_output_payload_state_index        (streamArbiter_20_io_output_payload_state_index    ), //o
    .io_output_payload_state_size         (streamArbiter_20_io_output_payload_state_size     ), //o
    .io_output_payload_state_id           (streamArbiter_20_io_output_payload_state_id       ), //o
    .io_output_payload_state_element      (streamArbiter_20_io_output_payload_state_element  ), //o
    .io_chosen                            (streamArbiter_20_io_chosen                        ), //o
    .io_chosenOH                          (streamArbiter_20_io_chosenOH                      ), //o
    .clk                                  (clk                                               ), //i
    .reset                                (reset                                             )  //i
  );
  assign inputs_0_valid = io_input_valid;
  assign inputs_0_payload_round_index = io_input_payload_round_index;
  assign inputs_0_payload_state_size = io_input_payload_state_size;
  assign inputs_0_payload_state_id = io_input_payload_state_id;
  assign inputs_0_payload_state_index = 4'b0000;
  assign inputs_0_payload_state_element = io_input_payload_state_elements_0;
  assign inputs_1_valid = io_input_valid;
  assign inputs_1_payload_round_index = io_input_payload_round_index;
  assign inputs_1_payload_state_size = io_input_payload_state_size;
  assign inputs_1_payload_state_id = io_input_payload_state_id;
  assign inputs_1_payload_state_index = 4'b0001;
  assign inputs_1_payload_state_element = io_input_payload_state_elements_1;
  assign inputs_2_valid = io_input_valid;
  assign inputs_2_payload_round_index = io_input_payload_round_index;
  assign inputs_2_payload_state_size = io_input_payload_state_size;
  assign inputs_2_payload_state_id = io_input_payload_state_id;
  assign inputs_2_payload_state_index = 4'b0010;
  assign inputs_2_payload_state_element = io_input_payload_state_elements_2;
  assign inputs_3_valid = io_input_valid;
  assign inputs_3_payload_round_index = io_input_payload_round_index;
  assign inputs_3_payload_state_size = io_input_payload_state_size;
  assign inputs_3_payload_state_id = io_input_payload_state_id;
  assign inputs_3_payload_state_index = 4'b0011;
  assign inputs_3_payload_state_element = io_input_payload_state_elements_3;
  assign inputs_4_valid = io_input_valid;
  assign inputs_4_payload_round_index = io_input_payload_round_index;
  assign inputs_4_payload_state_size = io_input_payload_state_size;
  assign inputs_4_payload_state_id = io_input_payload_state_id;
  assign inputs_4_payload_state_index = 4'b0100;
  assign inputs_4_payload_state_element = io_input_payload_state_elements_4;
  assign inputs_5_valid = io_input_valid;
  assign inputs_5_payload_round_index = io_input_payload_round_index;
  assign inputs_5_payload_state_size = io_input_payload_state_size;
  assign inputs_5_payload_state_id = io_input_payload_state_id;
  assign inputs_5_payload_state_index = 4'b0101;
  assign inputs_5_payload_state_element = io_input_payload_state_elements_5;
  assign inputs_6_valid = io_input_valid;
  assign inputs_6_payload_round_index = io_input_payload_round_index;
  assign inputs_6_payload_state_size = io_input_payload_state_size;
  assign inputs_6_payload_state_id = io_input_payload_state_id;
  assign inputs_6_payload_state_index = 4'b0110;
  assign inputs_6_payload_state_element = io_input_payload_state_elements_6;
  assign inputs_7_valid = io_input_valid;
  assign inputs_7_payload_round_index = io_input_payload_round_index;
  assign inputs_7_payload_state_size = io_input_payload_state_size;
  assign inputs_7_payload_state_id = io_input_payload_state_id;
  assign inputs_7_payload_state_index = 4'b0111;
  assign inputs_7_payload_state_element = io_input_payload_state_elements_7;
  assign inputs_8_valid = io_input_valid;
  assign inputs_8_payload_round_index = io_input_payload_round_index;
  assign inputs_8_payload_state_size = io_input_payload_state_size;
  assign inputs_8_payload_state_id = io_input_payload_state_id;
  assign inputs_8_payload_state_index = 4'b1000;
  assign inputs_8_payload_state_element = io_input_payload_state_elements_8;
  assign inputs_9_valid = io_input_valid;
  assign inputs_9_payload_round_index = io_input_payload_round_index;
  assign inputs_9_payload_state_size = io_input_payload_state_size;
  assign inputs_9_payload_state_id = io_input_payload_state_id;
  assign inputs_9_payload_state_index = 4'b1001;
  assign inputs_9_payload_state_element = io_input_payload_state_elements_9;
  assign inputs_10_valid = io_input_valid;
  assign inputs_10_payload_round_index = io_input_payload_round_index;
  assign inputs_10_payload_state_size = io_input_payload_state_size;
  assign inputs_10_payload_state_id = io_input_payload_state_id;
  assign inputs_10_payload_state_index = 4'b1010;
  assign inputs_10_payload_state_element = io_input_payload_state_elements_10;
  assign inputs_11_valid = io_input_valid;
  assign inputs_11_payload_round_index = io_input_payload_round_index;
  assign inputs_11_payload_state_size = io_input_payload_state_size;
  assign inputs_11_payload_state_id = io_input_payload_state_id;
  assign inputs_11_payload_state_index = 4'b1011;
  assign inputs_11_payload_state_element = io_input_payload_state_elements_11;
  assign io_input_ready = ({inputs_11_ready,{inputs_10_ready,{inputs_9_ready,{inputs_8_ready,{inputs_7_ready,{inputs_6_ready,{inputs_5_ready,{inputs_4_ready,{inputs_3_ready,{_zz_io_input_ready,_zz_io_input_ready_1}}}}}}}}}} == 12'hfff);
  always @(*) begin
    inputs_0_ready = inputs_0_m2sPipe_ready;
    if(when_Stream_l342) begin
      inputs_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! inputs_0_m2sPipe_valid);
  assign inputs_0_m2sPipe_valid = inputs_0_rValid;
  assign inputs_0_m2sPipe_payload_round_index = inputs_0_rData_round_index;
  assign inputs_0_m2sPipe_payload_state_index = inputs_0_rData_state_index;
  assign inputs_0_m2sPipe_payload_state_size = inputs_0_rData_state_size;
  assign inputs_0_m2sPipe_payload_state_id = inputs_0_rData_state_id;
  assign inputs_0_m2sPipe_payload_state_element = inputs_0_rData_state_element;
  assign buffer0_0_valid = inputs_0_m2sPipe_valid;
  assign inputs_0_m2sPipe_ready = buffer0_0_ready;
  assign buffer0_0_payload_round_index = inputs_0_m2sPipe_payload_round_index;
  assign buffer0_0_payload_state_index = inputs_0_m2sPipe_payload_state_index;
  assign buffer0_0_payload_state_size = inputs_0_m2sPipe_payload_state_size;
  assign buffer0_0_payload_state_id = inputs_0_m2sPipe_payload_state_id;
  assign buffer0_0_payload_state_element = inputs_0_m2sPipe_payload_state_element;
  assign when_Stream_l408 = (io_input_payload_state_size < 4'b0101);
  always @(*) begin
    inputs_3_thrown_valid = inputs_3_valid;
    if(when_Stream_l408) begin
      inputs_3_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_3_ready = inputs_3_thrown_ready;
    if(when_Stream_l408) begin
      inputs_3_ready = 1'b1;
    end
  end

  assign inputs_3_thrown_payload_round_index = inputs_3_payload_round_index;
  assign inputs_3_thrown_payload_state_index = inputs_3_payload_state_index;
  assign inputs_3_thrown_payload_state_size = inputs_3_payload_state_size;
  assign inputs_3_thrown_payload_state_id = inputs_3_payload_state_id;
  assign inputs_3_thrown_payload_state_element = inputs_3_payload_state_element;
  assign buffer0_0_ready = streamArbiter_12_io_inputs_0_ready;
  assign inputs_3_thrown_ready = streamArbiter_12_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_12_io_output_ready = streamArbiter_12_io_output_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      streamArbiter_12_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! streamArbiter_12_io_output_m2sPipe_valid);
  assign streamArbiter_12_io_output_m2sPipe_valid = streamArbiter_12_io_output_rValid;
  assign streamArbiter_12_io_output_m2sPipe_payload_round_index = streamArbiter_12_io_output_rData_round_index;
  assign streamArbiter_12_io_output_m2sPipe_payload_state_index = streamArbiter_12_io_output_rData_state_index;
  assign streamArbiter_12_io_output_m2sPipe_payload_state_size = streamArbiter_12_io_output_rData_state_size;
  assign streamArbiter_12_io_output_m2sPipe_payload_state_id = streamArbiter_12_io_output_rData_state_id;
  assign streamArbiter_12_io_output_m2sPipe_payload_state_element = streamArbiter_12_io_output_rData_state_element;
  assign buffer1_0_valid = streamArbiter_12_io_output_m2sPipe_valid;
  assign streamArbiter_12_io_output_m2sPipe_ready = buffer1_0_ready;
  assign buffer1_0_payload_round_index = streamArbiter_12_io_output_m2sPipe_payload_round_index;
  assign buffer1_0_payload_state_index = streamArbiter_12_io_output_m2sPipe_payload_state_index;
  assign buffer1_0_payload_state_size = streamArbiter_12_io_output_m2sPipe_payload_state_size;
  assign buffer1_0_payload_state_id = streamArbiter_12_io_output_m2sPipe_payload_state_id;
  assign buffer1_0_payload_state_element = streamArbiter_12_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_1 = (io_input_payload_state_size < 4'b1001);
  always @(*) begin
    inputs_6_thrown_valid = inputs_6_valid;
    if(when_Stream_l408_1) begin
      inputs_6_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_6_ready = inputs_6_thrown_ready;
    if(when_Stream_l408_1) begin
      inputs_6_ready = 1'b1;
    end
  end

  assign inputs_6_thrown_payload_round_index = inputs_6_payload_round_index;
  assign inputs_6_thrown_payload_state_index = inputs_6_payload_state_index;
  assign inputs_6_thrown_payload_state_size = inputs_6_payload_state_size;
  assign inputs_6_thrown_payload_state_id = inputs_6_payload_state_id;
  assign inputs_6_thrown_payload_state_element = inputs_6_payload_state_element;
  assign buffer1_0_ready = streamArbiter_13_io_inputs_0_ready;
  assign inputs_6_thrown_ready = streamArbiter_13_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_13_io_output_ready = streamArbiter_13_io_output_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      streamArbiter_13_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! streamArbiter_13_io_output_m2sPipe_valid);
  assign streamArbiter_13_io_output_m2sPipe_valid = streamArbiter_13_io_output_rValid;
  assign streamArbiter_13_io_output_m2sPipe_payload_round_index = streamArbiter_13_io_output_rData_round_index;
  assign streamArbiter_13_io_output_m2sPipe_payload_state_index = streamArbiter_13_io_output_rData_state_index;
  assign streamArbiter_13_io_output_m2sPipe_payload_state_size = streamArbiter_13_io_output_rData_state_size;
  assign streamArbiter_13_io_output_m2sPipe_payload_state_id = streamArbiter_13_io_output_rData_state_id;
  assign streamArbiter_13_io_output_m2sPipe_payload_state_element = streamArbiter_13_io_output_rData_state_element;
  assign buffer2_0_valid = streamArbiter_13_io_output_m2sPipe_valid;
  assign streamArbiter_13_io_output_m2sPipe_ready = buffer2_0_ready;
  assign buffer2_0_payload_round_index = streamArbiter_13_io_output_m2sPipe_payload_round_index;
  assign buffer2_0_payload_state_index = streamArbiter_13_io_output_m2sPipe_payload_state_index;
  assign buffer2_0_payload_state_size = streamArbiter_13_io_output_m2sPipe_payload_state_size;
  assign buffer2_0_payload_state_id = streamArbiter_13_io_output_m2sPipe_payload_state_id;
  assign buffer2_0_payload_state_element = streamArbiter_13_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_2 = (io_input_payload_state_size < 4'b1100);
  always @(*) begin
    inputs_9_thrown_valid = inputs_9_valid;
    if(when_Stream_l408_2) begin
      inputs_9_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_9_ready = inputs_9_thrown_ready;
    if(when_Stream_l408_2) begin
      inputs_9_ready = 1'b1;
    end
  end

  assign inputs_9_thrown_payload_round_index = inputs_9_payload_round_index;
  assign inputs_9_thrown_payload_state_index = inputs_9_payload_state_index;
  assign inputs_9_thrown_payload_state_size = inputs_9_payload_state_size;
  assign inputs_9_thrown_payload_state_id = inputs_9_payload_state_id;
  assign inputs_9_thrown_payload_state_element = inputs_9_payload_state_element;
  assign buffer2_0_ready = streamArbiter_14_io_inputs_0_ready;
  assign inputs_9_thrown_ready = streamArbiter_14_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_14_io_output_ready = streamArbiter_14_io_output_m2sPipe_ready;
    if(when_Stream_l342_3) begin
      streamArbiter_14_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! streamArbiter_14_io_output_m2sPipe_valid);
  assign streamArbiter_14_io_output_m2sPipe_valid = streamArbiter_14_io_output_rValid;
  assign streamArbiter_14_io_output_m2sPipe_payload_round_index = streamArbiter_14_io_output_rData_round_index;
  assign streamArbiter_14_io_output_m2sPipe_payload_state_index = streamArbiter_14_io_output_rData_state_index;
  assign streamArbiter_14_io_output_m2sPipe_payload_state_size = streamArbiter_14_io_output_rData_state_size;
  assign streamArbiter_14_io_output_m2sPipe_payload_state_id = streamArbiter_14_io_output_rData_state_id;
  assign streamArbiter_14_io_output_m2sPipe_payload_state_element = streamArbiter_14_io_output_rData_state_element;
  assign buffer3_0_valid = streamArbiter_14_io_output_m2sPipe_valid;
  assign streamArbiter_14_io_output_m2sPipe_ready = buffer3_0_ready;
  assign buffer3_0_payload_round_index = streamArbiter_14_io_output_m2sPipe_payload_round_index;
  assign buffer3_0_payload_state_index = streamArbiter_14_io_output_m2sPipe_payload_state_index;
  assign buffer3_0_payload_state_size = streamArbiter_14_io_output_m2sPipe_payload_state_size;
  assign buffer3_0_payload_state_id = streamArbiter_14_io_output_m2sPipe_payload_state_id;
  assign buffer3_0_payload_state_element = streamArbiter_14_io_output_m2sPipe_payload_state_element;
  always @(*) begin
    inputs_1_ready = inputs_1_m2sPipe_ready;
    if(when_Stream_l342_4) begin
      inputs_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_4 = (! inputs_1_m2sPipe_valid);
  assign inputs_1_m2sPipe_valid = inputs_1_rValid;
  assign inputs_1_m2sPipe_payload_round_index = inputs_1_rData_round_index;
  assign inputs_1_m2sPipe_payload_state_index = inputs_1_rData_state_index;
  assign inputs_1_m2sPipe_payload_state_size = inputs_1_rData_state_size;
  assign inputs_1_m2sPipe_payload_state_id = inputs_1_rData_state_id;
  assign inputs_1_m2sPipe_payload_state_element = inputs_1_rData_state_element;
  assign buffer0_1_valid = inputs_1_m2sPipe_valid;
  assign inputs_1_m2sPipe_ready = buffer0_1_ready;
  assign buffer0_1_payload_round_index = inputs_1_m2sPipe_payload_round_index;
  assign buffer0_1_payload_state_index = inputs_1_m2sPipe_payload_state_index;
  assign buffer0_1_payload_state_size = inputs_1_m2sPipe_payload_state_size;
  assign buffer0_1_payload_state_id = inputs_1_m2sPipe_payload_state_id;
  assign buffer0_1_payload_state_element = inputs_1_m2sPipe_payload_state_element;
  assign when_Stream_l408_3 = (io_input_payload_state_size < 4'b0101);
  always @(*) begin
    inputs_4_thrown_valid = inputs_4_valid;
    if(when_Stream_l408_3) begin
      inputs_4_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_4_ready = inputs_4_thrown_ready;
    if(when_Stream_l408_3) begin
      inputs_4_ready = 1'b1;
    end
  end

  assign inputs_4_thrown_payload_round_index = inputs_4_payload_round_index;
  assign inputs_4_thrown_payload_state_index = inputs_4_payload_state_index;
  assign inputs_4_thrown_payload_state_size = inputs_4_payload_state_size;
  assign inputs_4_thrown_payload_state_id = inputs_4_payload_state_id;
  assign inputs_4_thrown_payload_state_element = inputs_4_payload_state_element;
  assign buffer0_1_ready = streamArbiter_15_io_inputs_0_ready;
  assign inputs_4_thrown_ready = streamArbiter_15_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_15_io_output_ready = streamArbiter_15_io_output_m2sPipe_ready;
    if(when_Stream_l342_5) begin
      streamArbiter_15_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_5 = (! streamArbiter_15_io_output_m2sPipe_valid);
  assign streamArbiter_15_io_output_m2sPipe_valid = streamArbiter_15_io_output_rValid;
  assign streamArbiter_15_io_output_m2sPipe_payload_round_index = streamArbiter_15_io_output_rData_round_index;
  assign streamArbiter_15_io_output_m2sPipe_payload_state_index = streamArbiter_15_io_output_rData_state_index;
  assign streamArbiter_15_io_output_m2sPipe_payload_state_size = streamArbiter_15_io_output_rData_state_size;
  assign streamArbiter_15_io_output_m2sPipe_payload_state_id = streamArbiter_15_io_output_rData_state_id;
  assign streamArbiter_15_io_output_m2sPipe_payload_state_element = streamArbiter_15_io_output_rData_state_element;
  assign buffer1_1_valid = streamArbiter_15_io_output_m2sPipe_valid;
  assign streamArbiter_15_io_output_m2sPipe_ready = buffer1_1_ready;
  assign buffer1_1_payload_round_index = streamArbiter_15_io_output_m2sPipe_payload_round_index;
  assign buffer1_1_payload_state_index = streamArbiter_15_io_output_m2sPipe_payload_state_index;
  assign buffer1_1_payload_state_size = streamArbiter_15_io_output_m2sPipe_payload_state_size;
  assign buffer1_1_payload_state_id = streamArbiter_15_io_output_m2sPipe_payload_state_id;
  assign buffer1_1_payload_state_element = streamArbiter_15_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_4 = (io_input_payload_state_size < 4'b1001);
  always @(*) begin
    inputs_7_thrown_valid = inputs_7_valid;
    if(when_Stream_l408_4) begin
      inputs_7_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_7_ready = inputs_7_thrown_ready;
    if(when_Stream_l408_4) begin
      inputs_7_ready = 1'b1;
    end
  end

  assign inputs_7_thrown_payload_round_index = inputs_7_payload_round_index;
  assign inputs_7_thrown_payload_state_index = inputs_7_payload_state_index;
  assign inputs_7_thrown_payload_state_size = inputs_7_payload_state_size;
  assign inputs_7_thrown_payload_state_id = inputs_7_payload_state_id;
  assign inputs_7_thrown_payload_state_element = inputs_7_payload_state_element;
  assign buffer1_1_ready = streamArbiter_16_io_inputs_0_ready;
  assign inputs_7_thrown_ready = streamArbiter_16_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_16_io_output_ready = streamArbiter_16_io_output_m2sPipe_ready;
    if(when_Stream_l342_6) begin
      streamArbiter_16_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_6 = (! streamArbiter_16_io_output_m2sPipe_valid);
  assign streamArbiter_16_io_output_m2sPipe_valid = streamArbiter_16_io_output_rValid;
  assign streamArbiter_16_io_output_m2sPipe_payload_round_index = streamArbiter_16_io_output_rData_round_index;
  assign streamArbiter_16_io_output_m2sPipe_payload_state_index = streamArbiter_16_io_output_rData_state_index;
  assign streamArbiter_16_io_output_m2sPipe_payload_state_size = streamArbiter_16_io_output_rData_state_size;
  assign streamArbiter_16_io_output_m2sPipe_payload_state_id = streamArbiter_16_io_output_rData_state_id;
  assign streamArbiter_16_io_output_m2sPipe_payload_state_element = streamArbiter_16_io_output_rData_state_element;
  assign buffer2_1_valid = streamArbiter_16_io_output_m2sPipe_valid;
  assign streamArbiter_16_io_output_m2sPipe_ready = buffer2_1_ready;
  assign buffer2_1_payload_round_index = streamArbiter_16_io_output_m2sPipe_payload_round_index;
  assign buffer2_1_payload_state_index = streamArbiter_16_io_output_m2sPipe_payload_state_index;
  assign buffer2_1_payload_state_size = streamArbiter_16_io_output_m2sPipe_payload_state_size;
  assign buffer2_1_payload_state_id = streamArbiter_16_io_output_m2sPipe_payload_state_id;
  assign buffer2_1_payload_state_element = streamArbiter_16_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_5 = (io_input_payload_state_size < 4'b1100);
  always @(*) begin
    inputs_10_thrown_valid = inputs_10_valid;
    if(when_Stream_l408_5) begin
      inputs_10_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_10_ready = inputs_10_thrown_ready;
    if(when_Stream_l408_5) begin
      inputs_10_ready = 1'b1;
    end
  end

  assign inputs_10_thrown_payload_round_index = inputs_10_payload_round_index;
  assign inputs_10_thrown_payload_state_index = inputs_10_payload_state_index;
  assign inputs_10_thrown_payload_state_size = inputs_10_payload_state_size;
  assign inputs_10_thrown_payload_state_id = inputs_10_payload_state_id;
  assign inputs_10_thrown_payload_state_element = inputs_10_payload_state_element;
  assign buffer2_1_ready = streamArbiter_17_io_inputs_0_ready;
  assign inputs_10_thrown_ready = streamArbiter_17_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_17_io_output_ready = streamArbiter_17_io_output_m2sPipe_ready;
    if(when_Stream_l342_7) begin
      streamArbiter_17_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_7 = (! streamArbiter_17_io_output_m2sPipe_valid);
  assign streamArbiter_17_io_output_m2sPipe_valid = streamArbiter_17_io_output_rValid;
  assign streamArbiter_17_io_output_m2sPipe_payload_round_index = streamArbiter_17_io_output_rData_round_index;
  assign streamArbiter_17_io_output_m2sPipe_payload_state_index = streamArbiter_17_io_output_rData_state_index;
  assign streamArbiter_17_io_output_m2sPipe_payload_state_size = streamArbiter_17_io_output_rData_state_size;
  assign streamArbiter_17_io_output_m2sPipe_payload_state_id = streamArbiter_17_io_output_rData_state_id;
  assign streamArbiter_17_io_output_m2sPipe_payload_state_element = streamArbiter_17_io_output_rData_state_element;
  assign buffer3_1_valid = streamArbiter_17_io_output_m2sPipe_valid;
  assign streamArbiter_17_io_output_m2sPipe_ready = buffer3_1_ready;
  assign buffer3_1_payload_round_index = streamArbiter_17_io_output_m2sPipe_payload_round_index;
  assign buffer3_1_payload_state_index = streamArbiter_17_io_output_m2sPipe_payload_state_index;
  assign buffer3_1_payload_state_size = streamArbiter_17_io_output_m2sPipe_payload_state_size;
  assign buffer3_1_payload_state_id = streamArbiter_17_io_output_m2sPipe_payload_state_id;
  assign buffer3_1_payload_state_element = streamArbiter_17_io_output_m2sPipe_payload_state_element;
  always @(*) begin
    inputs_2_ready = inputs_2_m2sPipe_ready;
    if(when_Stream_l342_8) begin
      inputs_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_8 = (! inputs_2_m2sPipe_valid);
  assign inputs_2_m2sPipe_valid = inputs_2_rValid;
  assign inputs_2_m2sPipe_payload_round_index = inputs_2_rData_round_index;
  assign inputs_2_m2sPipe_payload_state_index = inputs_2_rData_state_index;
  assign inputs_2_m2sPipe_payload_state_size = inputs_2_rData_state_size;
  assign inputs_2_m2sPipe_payload_state_id = inputs_2_rData_state_id;
  assign inputs_2_m2sPipe_payload_state_element = inputs_2_rData_state_element;
  assign buffer0_2_valid = inputs_2_m2sPipe_valid;
  assign inputs_2_m2sPipe_ready = buffer0_2_ready;
  assign buffer0_2_payload_round_index = inputs_2_m2sPipe_payload_round_index;
  assign buffer0_2_payload_state_index = inputs_2_m2sPipe_payload_state_index;
  assign buffer0_2_payload_state_size = inputs_2_m2sPipe_payload_state_size;
  assign buffer0_2_payload_state_id = inputs_2_m2sPipe_payload_state_id;
  assign buffer0_2_payload_state_element = inputs_2_m2sPipe_payload_state_element;
  assign when_Stream_l408_6 = (io_input_payload_state_size < 4'b0101);
  always @(*) begin
    inputs_5_thrown_valid = inputs_5_valid;
    if(when_Stream_l408_6) begin
      inputs_5_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_5_ready = inputs_5_thrown_ready;
    if(when_Stream_l408_6) begin
      inputs_5_ready = 1'b1;
    end
  end

  assign inputs_5_thrown_payload_round_index = inputs_5_payload_round_index;
  assign inputs_5_thrown_payload_state_index = inputs_5_payload_state_index;
  assign inputs_5_thrown_payload_state_size = inputs_5_payload_state_size;
  assign inputs_5_thrown_payload_state_id = inputs_5_payload_state_id;
  assign inputs_5_thrown_payload_state_element = inputs_5_payload_state_element;
  assign buffer0_2_ready = streamArbiter_18_io_inputs_0_ready;
  assign inputs_5_thrown_ready = streamArbiter_18_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_18_io_output_ready = streamArbiter_18_io_output_m2sPipe_ready;
    if(when_Stream_l342_9) begin
      streamArbiter_18_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_9 = (! streamArbiter_18_io_output_m2sPipe_valid);
  assign streamArbiter_18_io_output_m2sPipe_valid = streamArbiter_18_io_output_rValid;
  assign streamArbiter_18_io_output_m2sPipe_payload_round_index = streamArbiter_18_io_output_rData_round_index;
  assign streamArbiter_18_io_output_m2sPipe_payload_state_index = streamArbiter_18_io_output_rData_state_index;
  assign streamArbiter_18_io_output_m2sPipe_payload_state_size = streamArbiter_18_io_output_rData_state_size;
  assign streamArbiter_18_io_output_m2sPipe_payload_state_id = streamArbiter_18_io_output_rData_state_id;
  assign streamArbiter_18_io_output_m2sPipe_payload_state_element = streamArbiter_18_io_output_rData_state_element;
  assign buffer1_2_valid = streamArbiter_18_io_output_m2sPipe_valid;
  assign streamArbiter_18_io_output_m2sPipe_ready = buffer1_2_ready;
  assign buffer1_2_payload_round_index = streamArbiter_18_io_output_m2sPipe_payload_round_index;
  assign buffer1_2_payload_state_index = streamArbiter_18_io_output_m2sPipe_payload_state_index;
  assign buffer1_2_payload_state_size = streamArbiter_18_io_output_m2sPipe_payload_state_size;
  assign buffer1_2_payload_state_id = streamArbiter_18_io_output_m2sPipe_payload_state_id;
  assign buffer1_2_payload_state_element = streamArbiter_18_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_7 = (io_input_payload_state_size < 4'b1001);
  always @(*) begin
    inputs_8_thrown_valid = inputs_8_valid;
    if(when_Stream_l408_7) begin
      inputs_8_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_8_ready = inputs_8_thrown_ready;
    if(when_Stream_l408_7) begin
      inputs_8_ready = 1'b1;
    end
  end

  assign inputs_8_thrown_payload_round_index = inputs_8_payload_round_index;
  assign inputs_8_thrown_payload_state_index = inputs_8_payload_state_index;
  assign inputs_8_thrown_payload_state_size = inputs_8_payload_state_size;
  assign inputs_8_thrown_payload_state_id = inputs_8_payload_state_id;
  assign inputs_8_thrown_payload_state_element = inputs_8_payload_state_element;
  assign buffer1_2_ready = streamArbiter_19_io_inputs_0_ready;
  assign inputs_8_thrown_ready = streamArbiter_19_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_19_io_output_ready = streamArbiter_19_io_output_m2sPipe_ready;
    if(when_Stream_l342_10) begin
      streamArbiter_19_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_10 = (! streamArbiter_19_io_output_m2sPipe_valid);
  assign streamArbiter_19_io_output_m2sPipe_valid = streamArbiter_19_io_output_rValid;
  assign streamArbiter_19_io_output_m2sPipe_payload_round_index = streamArbiter_19_io_output_rData_round_index;
  assign streamArbiter_19_io_output_m2sPipe_payload_state_index = streamArbiter_19_io_output_rData_state_index;
  assign streamArbiter_19_io_output_m2sPipe_payload_state_size = streamArbiter_19_io_output_rData_state_size;
  assign streamArbiter_19_io_output_m2sPipe_payload_state_id = streamArbiter_19_io_output_rData_state_id;
  assign streamArbiter_19_io_output_m2sPipe_payload_state_element = streamArbiter_19_io_output_rData_state_element;
  assign buffer2_2_valid = streamArbiter_19_io_output_m2sPipe_valid;
  assign streamArbiter_19_io_output_m2sPipe_ready = buffer2_2_ready;
  assign buffer2_2_payload_round_index = streamArbiter_19_io_output_m2sPipe_payload_round_index;
  assign buffer2_2_payload_state_index = streamArbiter_19_io_output_m2sPipe_payload_state_index;
  assign buffer2_2_payload_state_size = streamArbiter_19_io_output_m2sPipe_payload_state_size;
  assign buffer2_2_payload_state_id = streamArbiter_19_io_output_m2sPipe_payload_state_id;
  assign buffer2_2_payload_state_element = streamArbiter_19_io_output_m2sPipe_payload_state_element;
  assign when_Stream_l408_8 = (io_input_payload_state_size < 4'b1100);
  always @(*) begin
    inputs_11_thrown_valid = inputs_11_valid;
    if(when_Stream_l408_8) begin
      inputs_11_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    inputs_11_ready = inputs_11_thrown_ready;
    if(when_Stream_l408_8) begin
      inputs_11_ready = 1'b1;
    end
  end

  assign inputs_11_thrown_payload_round_index = inputs_11_payload_round_index;
  assign inputs_11_thrown_payload_state_index = inputs_11_payload_state_index;
  assign inputs_11_thrown_payload_state_size = inputs_11_payload_state_size;
  assign inputs_11_thrown_payload_state_id = inputs_11_payload_state_id;
  assign inputs_11_thrown_payload_state_element = inputs_11_payload_state_element;
  assign buffer2_2_ready = streamArbiter_20_io_inputs_0_ready;
  assign inputs_11_thrown_ready = streamArbiter_20_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_20_io_output_ready = streamArbiter_20_io_output_m2sPipe_ready;
    if(when_Stream_l342_11) begin
      streamArbiter_20_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_11 = (! streamArbiter_20_io_output_m2sPipe_valid);
  assign streamArbiter_20_io_output_m2sPipe_valid = streamArbiter_20_io_output_rValid;
  assign streamArbiter_20_io_output_m2sPipe_payload_round_index = streamArbiter_20_io_output_rData_round_index;
  assign streamArbiter_20_io_output_m2sPipe_payload_state_index = streamArbiter_20_io_output_rData_state_index;
  assign streamArbiter_20_io_output_m2sPipe_payload_state_size = streamArbiter_20_io_output_rData_state_size;
  assign streamArbiter_20_io_output_m2sPipe_payload_state_id = streamArbiter_20_io_output_rData_state_id;
  assign streamArbiter_20_io_output_m2sPipe_payload_state_element = streamArbiter_20_io_output_rData_state_element;
  assign buffer3_2_valid = streamArbiter_20_io_output_m2sPipe_valid;
  assign streamArbiter_20_io_output_m2sPipe_ready = buffer3_2_ready;
  assign buffer3_2_payload_round_index = streamArbiter_20_io_output_m2sPipe_payload_round_index;
  assign buffer3_2_payload_state_index = streamArbiter_20_io_output_m2sPipe_payload_state_index;
  assign buffer3_2_payload_state_size = streamArbiter_20_io_output_m2sPipe_payload_state_size;
  assign buffer3_2_payload_state_id = streamArbiter_20_io_output_m2sPipe_payload_state_id;
  assign buffer3_2_payload_state_element = streamArbiter_20_io_output_m2sPipe_payload_state_element;
  always @(*) begin
    buffer3_0_ready = buffer3_0_m2sPipe_ready;
    if(when_Stream_l342_12) begin
      buffer3_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_12 = (! buffer3_0_m2sPipe_valid);
  assign buffer3_0_m2sPipe_valid = buffer3_0_rValid;
  assign buffer3_0_m2sPipe_payload_round_index = buffer3_0_rData_round_index;
  assign buffer3_0_m2sPipe_payload_state_index = buffer3_0_rData_state_index;
  assign buffer3_0_m2sPipe_payload_state_size = buffer3_0_rData_state_size;
  assign buffer3_0_m2sPipe_payload_state_id = buffer3_0_rData_state_id;
  assign buffer3_0_m2sPipe_payload_state_element = buffer3_0_rData_state_element;
  assign buffers_0_0_valid = buffer3_0_m2sPipe_valid;
  assign buffer3_0_m2sPipe_ready = buffers_0_0_ready;
  assign buffers_0_0_payload_round_index = buffer3_0_m2sPipe_payload_round_index;
  assign buffers_0_0_payload_state_index = buffer3_0_m2sPipe_payload_state_index;
  assign buffers_0_0_payload_state_size = buffer3_0_m2sPipe_payload_state_size;
  assign buffers_0_0_payload_state_id = buffer3_0_m2sPipe_payload_state_id;
  assign buffers_0_0_payload_state_element = buffer3_0_m2sPipe_payload_state_element;
  always @(*) begin
    buffer3_1_ready = buffer3_1_m2sPipe_ready;
    if(when_Stream_l342_13) begin
      buffer3_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_13 = (! buffer3_1_m2sPipe_valid);
  assign buffer3_1_m2sPipe_valid = buffer3_1_rValid;
  assign buffer3_1_m2sPipe_payload_round_index = buffer3_1_rData_round_index;
  assign buffer3_1_m2sPipe_payload_state_index = buffer3_1_rData_state_index;
  assign buffer3_1_m2sPipe_payload_state_size = buffer3_1_rData_state_size;
  assign buffer3_1_m2sPipe_payload_state_id = buffer3_1_rData_state_id;
  assign buffer3_1_m2sPipe_payload_state_element = buffer3_1_rData_state_element;
  assign buffers_0_1_valid = buffer3_1_m2sPipe_valid;
  assign buffer3_1_m2sPipe_ready = buffers_0_1_ready;
  assign buffers_0_1_payload_round_index = buffer3_1_m2sPipe_payload_round_index;
  assign buffers_0_1_payload_state_index = buffer3_1_m2sPipe_payload_state_index;
  assign buffers_0_1_payload_state_size = buffer3_1_m2sPipe_payload_state_size;
  assign buffers_0_1_payload_state_id = buffer3_1_m2sPipe_payload_state_id;
  assign buffers_0_1_payload_state_element = buffer3_1_m2sPipe_payload_state_element;
  always @(*) begin
    buffer3_2_ready = buffer3_2_m2sPipe_ready;
    if(when_Stream_l342_14) begin
      buffer3_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_14 = (! buffer3_2_m2sPipe_valid);
  assign buffer3_2_m2sPipe_valid = buffer3_2_rValid;
  assign buffer3_2_m2sPipe_payload_round_index = buffer3_2_rData_round_index;
  assign buffer3_2_m2sPipe_payload_state_index = buffer3_2_rData_state_index;
  assign buffer3_2_m2sPipe_payload_state_size = buffer3_2_rData_state_size;
  assign buffer3_2_m2sPipe_payload_state_id = buffer3_2_rData_state_id;
  assign buffer3_2_m2sPipe_payload_state_element = buffer3_2_rData_state_element;
  assign buffers_0_2_valid = buffer3_2_m2sPipe_valid;
  assign buffer3_2_m2sPipe_ready = buffers_0_2_ready;
  assign buffers_0_2_payload_round_index = buffer3_2_m2sPipe_payload_round_index;
  assign buffers_0_2_payload_state_index = buffer3_2_m2sPipe_payload_state_index;
  assign buffers_0_2_payload_state_size = buffer3_2_m2sPipe_payload_state_size;
  assign buffers_0_2_payload_state_id = buffer3_2_m2sPipe_payload_state_id;
  assign buffers_0_2_payload_state_element = buffer3_2_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_0_0_ready = buffers_0_0_m2sPipe_ready;
    if(when_Stream_l342_15) begin
      buffers_0_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_15 = (! buffers_0_0_m2sPipe_valid);
  assign buffers_0_0_m2sPipe_valid = buffers_0_0_rValid;
  assign buffers_0_0_m2sPipe_payload_round_index = buffers_0_0_rData_round_index;
  assign buffers_0_0_m2sPipe_payload_state_index = buffers_0_0_rData_state_index;
  assign buffers_0_0_m2sPipe_payload_state_size = buffers_0_0_rData_state_size;
  assign buffers_0_0_m2sPipe_payload_state_id = buffers_0_0_rData_state_id;
  assign buffers_0_0_m2sPipe_payload_state_element = buffers_0_0_rData_state_element;
  assign buffers_1_0_valid = buffers_0_0_m2sPipe_valid;
  assign buffers_0_0_m2sPipe_ready = buffers_1_0_ready;
  assign buffers_1_0_payload_round_index = buffers_0_0_m2sPipe_payload_round_index;
  assign buffers_1_0_payload_state_index = buffers_0_0_m2sPipe_payload_state_index;
  assign buffers_1_0_payload_state_size = buffers_0_0_m2sPipe_payload_state_size;
  assign buffers_1_0_payload_state_id = buffers_0_0_m2sPipe_payload_state_id;
  assign buffers_1_0_payload_state_element = buffers_0_0_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_0_1_ready = buffers_0_1_m2sPipe_ready;
    if(when_Stream_l342_16) begin
      buffers_0_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_16 = (! buffers_0_1_m2sPipe_valid);
  assign buffers_0_1_m2sPipe_valid = buffers_0_1_rValid;
  assign buffers_0_1_m2sPipe_payload_round_index = buffers_0_1_rData_round_index;
  assign buffers_0_1_m2sPipe_payload_state_index = buffers_0_1_rData_state_index;
  assign buffers_0_1_m2sPipe_payload_state_size = buffers_0_1_rData_state_size;
  assign buffers_0_1_m2sPipe_payload_state_id = buffers_0_1_rData_state_id;
  assign buffers_0_1_m2sPipe_payload_state_element = buffers_0_1_rData_state_element;
  assign buffers_1_1_valid = buffers_0_1_m2sPipe_valid;
  assign buffers_0_1_m2sPipe_ready = buffers_1_1_ready;
  assign buffers_1_1_payload_round_index = buffers_0_1_m2sPipe_payload_round_index;
  assign buffers_1_1_payload_state_index = buffers_0_1_m2sPipe_payload_state_index;
  assign buffers_1_1_payload_state_size = buffers_0_1_m2sPipe_payload_state_size;
  assign buffers_1_1_payload_state_id = buffers_0_1_m2sPipe_payload_state_id;
  assign buffers_1_1_payload_state_element = buffers_0_1_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_0_2_ready = buffers_0_2_m2sPipe_ready;
    if(when_Stream_l342_17) begin
      buffers_0_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_17 = (! buffers_0_2_m2sPipe_valid);
  assign buffers_0_2_m2sPipe_valid = buffers_0_2_rValid;
  assign buffers_0_2_m2sPipe_payload_round_index = buffers_0_2_rData_round_index;
  assign buffers_0_2_m2sPipe_payload_state_index = buffers_0_2_rData_state_index;
  assign buffers_0_2_m2sPipe_payload_state_size = buffers_0_2_rData_state_size;
  assign buffers_0_2_m2sPipe_payload_state_id = buffers_0_2_rData_state_id;
  assign buffers_0_2_m2sPipe_payload_state_element = buffers_0_2_rData_state_element;
  assign buffers_1_2_valid = buffers_0_2_m2sPipe_valid;
  assign buffers_0_2_m2sPipe_ready = buffers_1_2_ready;
  assign buffers_1_2_payload_round_index = buffers_0_2_m2sPipe_payload_round_index;
  assign buffers_1_2_payload_state_index = buffers_0_2_m2sPipe_payload_state_index;
  assign buffers_1_2_payload_state_size = buffers_0_2_m2sPipe_payload_state_size;
  assign buffers_1_2_payload_state_id = buffers_0_2_m2sPipe_payload_state_id;
  assign buffers_1_2_payload_state_element = buffers_0_2_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_1_0_ready = buffers_1_0_m2sPipe_ready;
    if(when_Stream_l342_18) begin
      buffers_1_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_18 = (! buffers_1_0_m2sPipe_valid);
  assign buffers_1_0_m2sPipe_valid = buffers_1_0_rValid;
  assign buffers_1_0_m2sPipe_payload_round_index = buffers_1_0_rData_round_index;
  assign buffers_1_0_m2sPipe_payload_state_index = buffers_1_0_rData_state_index;
  assign buffers_1_0_m2sPipe_payload_state_size = buffers_1_0_rData_state_size;
  assign buffers_1_0_m2sPipe_payload_state_id = buffers_1_0_rData_state_id;
  assign buffers_1_0_m2sPipe_payload_state_element = buffers_1_0_rData_state_element;
  assign buffers_2_0_valid = buffers_1_0_m2sPipe_valid;
  assign buffers_1_0_m2sPipe_ready = buffers_2_0_ready;
  assign buffers_2_0_payload_round_index = buffers_1_0_m2sPipe_payload_round_index;
  assign buffers_2_0_payload_state_index = buffers_1_0_m2sPipe_payload_state_index;
  assign buffers_2_0_payload_state_size = buffers_1_0_m2sPipe_payload_state_size;
  assign buffers_2_0_payload_state_id = buffers_1_0_m2sPipe_payload_state_id;
  assign buffers_2_0_payload_state_element = buffers_1_0_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_1_1_ready = buffers_1_1_m2sPipe_ready;
    if(when_Stream_l342_19) begin
      buffers_1_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_19 = (! buffers_1_1_m2sPipe_valid);
  assign buffers_1_1_m2sPipe_valid = buffers_1_1_rValid;
  assign buffers_1_1_m2sPipe_payload_round_index = buffers_1_1_rData_round_index;
  assign buffers_1_1_m2sPipe_payload_state_index = buffers_1_1_rData_state_index;
  assign buffers_1_1_m2sPipe_payload_state_size = buffers_1_1_rData_state_size;
  assign buffers_1_1_m2sPipe_payload_state_id = buffers_1_1_rData_state_id;
  assign buffers_1_1_m2sPipe_payload_state_element = buffers_1_1_rData_state_element;
  assign buffers_2_1_valid = buffers_1_1_m2sPipe_valid;
  assign buffers_1_1_m2sPipe_ready = buffers_2_1_ready;
  assign buffers_2_1_payload_round_index = buffers_1_1_m2sPipe_payload_round_index;
  assign buffers_2_1_payload_state_index = buffers_1_1_m2sPipe_payload_state_index;
  assign buffers_2_1_payload_state_size = buffers_1_1_m2sPipe_payload_state_size;
  assign buffers_2_1_payload_state_id = buffers_1_1_m2sPipe_payload_state_id;
  assign buffers_2_1_payload_state_element = buffers_1_1_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_1_2_ready = buffers_1_2_m2sPipe_ready;
    if(when_Stream_l342_20) begin
      buffers_1_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_20 = (! buffers_1_2_m2sPipe_valid);
  assign buffers_1_2_m2sPipe_valid = buffers_1_2_rValid;
  assign buffers_1_2_m2sPipe_payload_round_index = buffers_1_2_rData_round_index;
  assign buffers_1_2_m2sPipe_payload_state_index = buffers_1_2_rData_state_index;
  assign buffers_1_2_m2sPipe_payload_state_size = buffers_1_2_rData_state_size;
  assign buffers_1_2_m2sPipe_payload_state_id = buffers_1_2_rData_state_id;
  assign buffers_1_2_m2sPipe_payload_state_element = buffers_1_2_rData_state_element;
  assign buffers_2_2_valid = buffers_1_2_m2sPipe_valid;
  assign buffers_1_2_m2sPipe_ready = buffers_2_2_ready;
  assign buffers_2_2_payload_round_index = buffers_1_2_m2sPipe_payload_round_index;
  assign buffers_2_2_payload_state_index = buffers_1_2_m2sPipe_payload_state_index;
  assign buffers_2_2_payload_state_size = buffers_1_2_m2sPipe_payload_state_size;
  assign buffers_2_2_payload_state_id = buffers_1_2_m2sPipe_payload_state_id;
  assign buffers_2_2_payload_state_element = buffers_1_2_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_2_0_ready = buffers_2_0_m2sPipe_ready;
    if(when_Stream_l342_21) begin
      buffers_2_0_ready = 1'b1;
    end
  end

  assign when_Stream_l342_21 = (! buffers_2_0_m2sPipe_valid);
  assign buffers_2_0_m2sPipe_valid = buffers_2_0_rValid;
  assign buffers_2_0_m2sPipe_payload_round_index = buffers_2_0_rData_round_index;
  assign buffers_2_0_m2sPipe_payload_state_index = buffers_2_0_rData_state_index;
  assign buffers_2_0_m2sPipe_payload_state_size = buffers_2_0_rData_state_size;
  assign buffers_2_0_m2sPipe_payload_state_id = buffers_2_0_rData_state_id;
  assign buffers_2_0_m2sPipe_payload_state_element = buffers_2_0_rData_state_element;
  assign buffers_3_0_valid = buffers_2_0_m2sPipe_valid;
  assign buffers_2_0_m2sPipe_ready = buffers_3_0_ready;
  assign buffers_3_0_payload_round_index = buffers_2_0_m2sPipe_payload_round_index;
  assign buffers_3_0_payload_state_index = buffers_2_0_m2sPipe_payload_state_index;
  assign buffers_3_0_payload_state_size = buffers_2_0_m2sPipe_payload_state_size;
  assign buffers_3_0_payload_state_id = buffers_2_0_m2sPipe_payload_state_id;
  assign buffers_3_0_payload_state_element = buffers_2_0_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_2_1_ready = buffers_2_1_m2sPipe_ready;
    if(when_Stream_l342_22) begin
      buffers_2_1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_22 = (! buffers_2_1_m2sPipe_valid);
  assign buffers_2_1_m2sPipe_valid = buffers_2_1_rValid;
  assign buffers_2_1_m2sPipe_payload_round_index = buffers_2_1_rData_round_index;
  assign buffers_2_1_m2sPipe_payload_state_index = buffers_2_1_rData_state_index;
  assign buffers_2_1_m2sPipe_payload_state_size = buffers_2_1_rData_state_size;
  assign buffers_2_1_m2sPipe_payload_state_id = buffers_2_1_rData_state_id;
  assign buffers_2_1_m2sPipe_payload_state_element = buffers_2_1_rData_state_element;
  assign buffers_3_1_valid = buffers_2_1_m2sPipe_valid;
  assign buffers_2_1_m2sPipe_ready = buffers_3_1_ready;
  assign buffers_3_1_payload_round_index = buffers_2_1_m2sPipe_payload_round_index;
  assign buffers_3_1_payload_state_index = buffers_2_1_m2sPipe_payload_state_index;
  assign buffers_3_1_payload_state_size = buffers_2_1_m2sPipe_payload_state_size;
  assign buffers_3_1_payload_state_id = buffers_2_1_m2sPipe_payload_state_id;
  assign buffers_3_1_payload_state_element = buffers_2_1_m2sPipe_payload_state_element;
  always @(*) begin
    buffers_2_2_ready = buffers_2_2_m2sPipe_ready;
    if(when_Stream_l342_23) begin
      buffers_2_2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_23 = (! buffers_2_2_m2sPipe_valid);
  assign buffers_2_2_m2sPipe_valid = buffers_2_2_rValid;
  assign buffers_2_2_m2sPipe_payload_round_index = buffers_2_2_rData_round_index;
  assign buffers_2_2_m2sPipe_payload_state_index = buffers_2_2_rData_state_index;
  assign buffers_2_2_m2sPipe_payload_state_size = buffers_2_2_rData_state_size;
  assign buffers_2_2_m2sPipe_payload_state_id = buffers_2_2_rData_state_id;
  assign buffers_2_2_m2sPipe_payload_state_element = buffers_2_2_rData_state_element;
  assign buffers_3_2_valid = buffers_2_2_m2sPipe_valid;
  assign buffers_2_2_m2sPipe_ready = buffers_3_2_ready;
  assign buffers_3_2_payload_round_index = buffers_2_2_m2sPipe_payload_round_index;
  assign buffers_3_2_payload_state_index = buffers_2_2_m2sPipe_payload_state_index;
  assign buffers_3_2_payload_state_size = buffers_2_2_m2sPipe_payload_state_size;
  assign buffers_3_2_payload_state_id = buffers_2_2_m2sPipe_payload_state_id;
  assign buffers_3_2_payload_state_element = buffers_2_2_m2sPipe_payload_state_element;
  always @(*) begin
    io_residue = 4'b1100;
    if(when_PoseidonTopLevel_l90) begin
      io_residue = 4'b1001;
    end
    if(when_PoseidonTopLevel_l93) begin
      io_residue = 4'b0110;
    end
    if(when_PoseidonTopLevel_l96) begin
      io_residue = 4'b0011;
    end
    if(when_PoseidonTopLevel_l99) begin
      io_residue = 4'b0000;
    end
  end

  assign when_PoseidonTopLevel_l90 = ((buffers_0_0_valid && buffers_0_1_valid) && buffers_0_2_valid);
  assign when_PoseidonTopLevel_l93 = ((buffers_1_0_valid && buffers_1_1_valid) && buffers_1_2_valid);
  assign when_PoseidonTopLevel_l96 = ((buffers_2_0_valid && buffers_2_1_valid) && buffers_2_2_valid);
  assign when_PoseidonTopLevel_l99 = ((buffers_3_0_valid && buffers_3_1_valid) && buffers_3_2_valid);
  assign io_outputs_0_valid = buffers_3_0_valid;
  assign buffers_3_0_ready = io_outputs_0_ready;
  assign io_outputs_0_payload_round_index = buffers_3_0_payload_round_index;
  assign io_outputs_0_payload_state_index = buffers_3_0_payload_state_index;
  assign io_outputs_0_payload_state_size = buffers_3_0_payload_state_size;
  assign io_outputs_0_payload_state_id = buffers_3_0_payload_state_id;
  assign io_outputs_0_payload_state_element = buffers_3_0_payload_state_element;
  assign io_outputs_1_valid = buffers_3_1_valid;
  assign buffers_3_1_ready = io_outputs_1_ready;
  assign io_outputs_1_payload_round_index = buffers_3_1_payload_round_index;
  assign io_outputs_1_payload_state_index = buffers_3_1_payload_state_index;
  assign io_outputs_1_payload_state_size = buffers_3_1_payload_state_size;
  assign io_outputs_1_payload_state_id = buffers_3_1_payload_state_id;
  assign io_outputs_1_payload_state_element = buffers_3_1_payload_state_element;
  assign io_outputs_2_valid = buffers_3_2_valid;
  assign buffers_3_2_ready = io_outputs_2_ready;
  assign io_outputs_2_payload_round_index = buffers_3_2_payload_round_index;
  assign io_outputs_2_payload_state_index = buffers_3_2_payload_state_index;
  assign io_outputs_2_payload_state_size = buffers_3_2_payload_state_size;
  assign io_outputs_2_payload_state_id = buffers_3_2_payload_state_id;
  assign io_outputs_2_payload_state_element = buffers_3_2_payload_state_element;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      inputs_0_rValid <= 1'b0;
      streamArbiter_12_io_output_rValid <= 1'b0;
      streamArbiter_13_io_output_rValid <= 1'b0;
      streamArbiter_14_io_output_rValid <= 1'b0;
      inputs_1_rValid <= 1'b0;
      streamArbiter_15_io_output_rValid <= 1'b0;
      streamArbiter_16_io_output_rValid <= 1'b0;
      streamArbiter_17_io_output_rValid <= 1'b0;
      inputs_2_rValid <= 1'b0;
      streamArbiter_18_io_output_rValid <= 1'b0;
      streamArbiter_19_io_output_rValid <= 1'b0;
      streamArbiter_20_io_output_rValid <= 1'b0;
      buffer3_0_rValid <= 1'b0;
      buffer3_1_rValid <= 1'b0;
      buffer3_2_rValid <= 1'b0;
      buffers_0_0_rValid <= 1'b0;
      buffers_0_1_rValid <= 1'b0;
      buffers_0_2_rValid <= 1'b0;
      buffers_1_0_rValid <= 1'b0;
      buffers_1_1_rValid <= 1'b0;
      buffers_1_2_rValid <= 1'b0;
      buffers_2_0_rValid <= 1'b0;
      buffers_2_1_rValid <= 1'b0;
      buffers_2_2_rValid <= 1'b0;
    end else begin
      if(inputs_0_ready) begin
        inputs_0_rValid <= inputs_0_valid;
      end
      if(streamArbiter_12_io_output_ready) begin
        streamArbiter_12_io_output_rValid <= streamArbiter_12_io_output_valid;
      end
      if(streamArbiter_13_io_output_ready) begin
        streamArbiter_13_io_output_rValid <= streamArbiter_13_io_output_valid;
      end
      if(streamArbiter_14_io_output_ready) begin
        streamArbiter_14_io_output_rValid <= streamArbiter_14_io_output_valid;
      end
      if(inputs_1_ready) begin
        inputs_1_rValid <= inputs_1_valid;
      end
      if(streamArbiter_15_io_output_ready) begin
        streamArbiter_15_io_output_rValid <= streamArbiter_15_io_output_valid;
      end
      if(streamArbiter_16_io_output_ready) begin
        streamArbiter_16_io_output_rValid <= streamArbiter_16_io_output_valid;
      end
      if(streamArbiter_17_io_output_ready) begin
        streamArbiter_17_io_output_rValid <= streamArbiter_17_io_output_valid;
      end
      if(inputs_2_ready) begin
        inputs_2_rValid <= inputs_2_valid;
      end
      if(streamArbiter_18_io_output_ready) begin
        streamArbiter_18_io_output_rValid <= streamArbiter_18_io_output_valid;
      end
      if(streamArbiter_19_io_output_ready) begin
        streamArbiter_19_io_output_rValid <= streamArbiter_19_io_output_valid;
      end
      if(streamArbiter_20_io_output_ready) begin
        streamArbiter_20_io_output_rValid <= streamArbiter_20_io_output_valid;
      end
      if(buffer3_0_ready) begin
        buffer3_0_rValid <= buffer3_0_valid;
      end
      if(buffer3_1_ready) begin
        buffer3_1_rValid <= buffer3_1_valid;
      end
      if(buffer3_2_ready) begin
        buffer3_2_rValid <= buffer3_2_valid;
      end
      if(buffers_0_0_ready) begin
        buffers_0_0_rValid <= buffers_0_0_valid;
      end
      if(buffers_0_1_ready) begin
        buffers_0_1_rValid <= buffers_0_1_valid;
      end
      if(buffers_0_2_ready) begin
        buffers_0_2_rValid <= buffers_0_2_valid;
      end
      if(buffers_1_0_ready) begin
        buffers_1_0_rValid <= buffers_1_0_valid;
      end
      if(buffers_1_1_ready) begin
        buffers_1_1_rValid <= buffers_1_1_valid;
      end
      if(buffers_1_2_ready) begin
        buffers_1_2_rValid <= buffers_1_2_valid;
      end
      if(buffers_2_0_ready) begin
        buffers_2_0_rValid <= buffers_2_0_valid;
      end
      if(buffers_2_1_ready) begin
        buffers_2_1_rValid <= buffers_2_1_valid;
      end
      if(buffers_2_2_ready) begin
        buffers_2_2_rValid <= buffers_2_2_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(inputs_0_ready) begin
      inputs_0_rData_round_index <= inputs_0_payload_round_index;
      inputs_0_rData_state_index <= inputs_0_payload_state_index;
      inputs_0_rData_state_size <= inputs_0_payload_state_size;
      inputs_0_rData_state_id <= inputs_0_payload_state_id;
      inputs_0_rData_state_element <= inputs_0_payload_state_element;
    end
    if(streamArbiter_12_io_output_ready) begin
      streamArbiter_12_io_output_rData_round_index <= streamArbiter_12_io_output_payload_round_index;
      streamArbiter_12_io_output_rData_state_index <= streamArbiter_12_io_output_payload_state_index;
      streamArbiter_12_io_output_rData_state_size <= streamArbiter_12_io_output_payload_state_size;
      streamArbiter_12_io_output_rData_state_id <= streamArbiter_12_io_output_payload_state_id;
      streamArbiter_12_io_output_rData_state_element <= streamArbiter_12_io_output_payload_state_element;
    end
    if(streamArbiter_13_io_output_ready) begin
      streamArbiter_13_io_output_rData_round_index <= streamArbiter_13_io_output_payload_round_index;
      streamArbiter_13_io_output_rData_state_index <= streamArbiter_13_io_output_payload_state_index;
      streamArbiter_13_io_output_rData_state_size <= streamArbiter_13_io_output_payload_state_size;
      streamArbiter_13_io_output_rData_state_id <= streamArbiter_13_io_output_payload_state_id;
      streamArbiter_13_io_output_rData_state_element <= streamArbiter_13_io_output_payload_state_element;
    end
    if(streamArbiter_14_io_output_ready) begin
      streamArbiter_14_io_output_rData_round_index <= streamArbiter_14_io_output_payload_round_index;
      streamArbiter_14_io_output_rData_state_index <= streamArbiter_14_io_output_payload_state_index;
      streamArbiter_14_io_output_rData_state_size <= streamArbiter_14_io_output_payload_state_size;
      streamArbiter_14_io_output_rData_state_id <= streamArbiter_14_io_output_payload_state_id;
      streamArbiter_14_io_output_rData_state_element <= streamArbiter_14_io_output_payload_state_element;
    end
    if(inputs_1_ready) begin
      inputs_1_rData_round_index <= inputs_1_payload_round_index;
      inputs_1_rData_state_index <= inputs_1_payload_state_index;
      inputs_1_rData_state_size <= inputs_1_payload_state_size;
      inputs_1_rData_state_id <= inputs_1_payload_state_id;
      inputs_1_rData_state_element <= inputs_1_payload_state_element;
    end
    if(streamArbiter_15_io_output_ready) begin
      streamArbiter_15_io_output_rData_round_index <= streamArbiter_15_io_output_payload_round_index;
      streamArbiter_15_io_output_rData_state_index <= streamArbiter_15_io_output_payload_state_index;
      streamArbiter_15_io_output_rData_state_size <= streamArbiter_15_io_output_payload_state_size;
      streamArbiter_15_io_output_rData_state_id <= streamArbiter_15_io_output_payload_state_id;
      streamArbiter_15_io_output_rData_state_element <= streamArbiter_15_io_output_payload_state_element;
    end
    if(streamArbiter_16_io_output_ready) begin
      streamArbiter_16_io_output_rData_round_index <= streamArbiter_16_io_output_payload_round_index;
      streamArbiter_16_io_output_rData_state_index <= streamArbiter_16_io_output_payload_state_index;
      streamArbiter_16_io_output_rData_state_size <= streamArbiter_16_io_output_payload_state_size;
      streamArbiter_16_io_output_rData_state_id <= streamArbiter_16_io_output_payload_state_id;
      streamArbiter_16_io_output_rData_state_element <= streamArbiter_16_io_output_payload_state_element;
    end
    if(streamArbiter_17_io_output_ready) begin
      streamArbiter_17_io_output_rData_round_index <= streamArbiter_17_io_output_payload_round_index;
      streamArbiter_17_io_output_rData_state_index <= streamArbiter_17_io_output_payload_state_index;
      streamArbiter_17_io_output_rData_state_size <= streamArbiter_17_io_output_payload_state_size;
      streamArbiter_17_io_output_rData_state_id <= streamArbiter_17_io_output_payload_state_id;
      streamArbiter_17_io_output_rData_state_element <= streamArbiter_17_io_output_payload_state_element;
    end
    if(inputs_2_ready) begin
      inputs_2_rData_round_index <= inputs_2_payload_round_index;
      inputs_2_rData_state_index <= inputs_2_payload_state_index;
      inputs_2_rData_state_size <= inputs_2_payload_state_size;
      inputs_2_rData_state_id <= inputs_2_payload_state_id;
      inputs_2_rData_state_element <= inputs_2_payload_state_element;
    end
    if(streamArbiter_18_io_output_ready) begin
      streamArbiter_18_io_output_rData_round_index <= streamArbiter_18_io_output_payload_round_index;
      streamArbiter_18_io_output_rData_state_index <= streamArbiter_18_io_output_payload_state_index;
      streamArbiter_18_io_output_rData_state_size <= streamArbiter_18_io_output_payload_state_size;
      streamArbiter_18_io_output_rData_state_id <= streamArbiter_18_io_output_payload_state_id;
      streamArbiter_18_io_output_rData_state_element <= streamArbiter_18_io_output_payload_state_element;
    end
    if(streamArbiter_19_io_output_ready) begin
      streamArbiter_19_io_output_rData_round_index <= streamArbiter_19_io_output_payload_round_index;
      streamArbiter_19_io_output_rData_state_index <= streamArbiter_19_io_output_payload_state_index;
      streamArbiter_19_io_output_rData_state_size <= streamArbiter_19_io_output_payload_state_size;
      streamArbiter_19_io_output_rData_state_id <= streamArbiter_19_io_output_payload_state_id;
      streamArbiter_19_io_output_rData_state_element <= streamArbiter_19_io_output_payload_state_element;
    end
    if(streamArbiter_20_io_output_ready) begin
      streamArbiter_20_io_output_rData_round_index <= streamArbiter_20_io_output_payload_round_index;
      streamArbiter_20_io_output_rData_state_index <= streamArbiter_20_io_output_payload_state_index;
      streamArbiter_20_io_output_rData_state_size <= streamArbiter_20_io_output_payload_state_size;
      streamArbiter_20_io_output_rData_state_id <= streamArbiter_20_io_output_payload_state_id;
      streamArbiter_20_io_output_rData_state_element <= streamArbiter_20_io_output_payload_state_element;
    end
    if(buffer3_0_ready) begin
      buffer3_0_rData_round_index <= buffer3_0_payload_round_index;
      buffer3_0_rData_state_index <= buffer3_0_payload_state_index;
      buffer3_0_rData_state_size <= buffer3_0_payload_state_size;
      buffer3_0_rData_state_id <= buffer3_0_payload_state_id;
      buffer3_0_rData_state_element <= buffer3_0_payload_state_element;
    end
    if(buffer3_1_ready) begin
      buffer3_1_rData_round_index <= buffer3_1_payload_round_index;
      buffer3_1_rData_state_index <= buffer3_1_payload_state_index;
      buffer3_1_rData_state_size <= buffer3_1_payload_state_size;
      buffer3_1_rData_state_id <= buffer3_1_payload_state_id;
      buffer3_1_rData_state_element <= buffer3_1_payload_state_element;
    end
    if(buffer3_2_ready) begin
      buffer3_2_rData_round_index <= buffer3_2_payload_round_index;
      buffer3_2_rData_state_index <= buffer3_2_payload_state_index;
      buffer3_2_rData_state_size <= buffer3_2_payload_state_size;
      buffer3_2_rData_state_id <= buffer3_2_payload_state_id;
      buffer3_2_rData_state_element <= buffer3_2_payload_state_element;
    end
    if(buffers_0_0_ready) begin
      buffers_0_0_rData_round_index <= buffers_0_0_payload_round_index;
      buffers_0_0_rData_state_index <= buffers_0_0_payload_state_index;
      buffers_0_0_rData_state_size <= buffers_0_0_payload_state_size;
      buffers_0_0_rData_state_id <= buffers_0_0_payload_state_id;
      buffers_0_0_rData_state_element <= buffers_0_0_payload_state_element;
    end
    if(buffers_0_1_ready) begin
      buffers_0_1_rData_round_index <= buffers_0_1_payload_round_index;
      buffers_0_1_rData_state_index <= buffers_0_1_payload_state_index;
      buffers_0_1_rData_state_size <= buffers_0_1_payload_state_size;
      buffers_0_1_rData_state_id <= buffers_0_1_payload_state_id;
      buffers_0_1_rData_state_element <= buffers_0_1_payload_state_element;
    end
    if(buffers_0_2_ready) begin
      buffers_0_2_rData_round_index <= buffers_0_2_payload_round_index;
      buffers_0_2_rData_state_index <= buffers_0_2_payload_state_index;
      buffers_0_2_rData_state_size <= buffers_0_2_payload_state_size;
      buffers_0_2_rData_state_id <= buffers_0_2_payload_state_id;
      buffers_0_2_rData_state_element <= buffers_0_2_payload_state_element;
    end
    if(buffers_1_0_ready) begin
      buffers_1_0_rData_round_index <= buffers_1_0_payload_round_index;
      buffers_1_0_rData_state_index <= buffers_1_0_payload_state_index;
      buffers_1_0_rData_state_size <= buffers_1_0_payload_state_size;
      buffers_1_0_rData_state_id <= buffers_1_0_payload_state_id;
      buffers_1_0_rData_state_element <= buffers_1_0_payload_state_element;
    end
    if(buffers_1_1_ready) begin
      buffers_1_1_rData_round_index <= buffers_1_1_payload_round_index;
      buffers_1_1_rData_state_index <= buffers_1_1_payload_state_index;
      buffers_1_1_rData_state_size <= buffers_1_1_payload_state_size;
      buffers_1_1_rData_state_id <= buffers_1_1_payload_state_id;
      buffers_1_1_rData_state_element <= buffers_1_1_payload_state_element;
    end
    if(buffers_1_2_ready) begin
      buffers_1_2_rData_round_index <= buffers_1_2_payload_round_index;
      buffers_1_2_rData_state_index <= buffers_1_2_payload_state_index;
      buffers_1_2_rData_state_size <= buffers_1_2_payload_state_size;
      buffers_1_2_rData_state_id <= buffers_1_2_payload_state_id;
      buffers_1_2_rData_state_element <= buffers_1_2_payload_state_element;
    end
    if(buffers_2_0_ready) begin
      buffers_2_0_rData_round_index <= buffers_2_0_payload_round_index;
      buffers_2_0_rData_state_index <= buffers_2_0_payload_state_index;
      buffers_2_0_rData_state_size <= buffers_2_0_payload_state_size;
      buffers_2_0_rData_state_id <= buffers_2_0_payload_state_id;
      buffers_2_0_rData_state_element <= buffers_2_0_payload_state_element;
    end
    if(buffers_2_1_ready) begin
      buffers_2_1_rData_round_index <= buffers_2_1_payload_round_index;
      buffers_2_1_rData_state_index <= buffers_2_1_payload_state_index;
      buffers_2_1_rData_state_size <= buffers_2_1_payload_state_size;
      buffers_2_1_rData_state_id <= buffers_2_1_payload_state_id;
      buffers_2_1_rData_state_element <= buffers_2_1_payload_state_element;
    end
    if(buffers_2_2_ready) begin
      buffers_2_2_rData_round_index <= buffers_2_2_payload_round_index;
      buffers_2_2_rData_state_index <= buffers_2_2_payload_state_index;
      buffers_2_2_rData_state_size <= buffers_2_2_payload_state_size;
      buffers_2_2_rData_state_id <= buffers_2_2_payload_state_id;
      buffers_2_2_rData_state_element <= buffers_2_2_payload_state_element;
    end
  end


endmodule

module PoseidonThread_2 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index;
  wire       [2:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index;
  reg        [254:0]  AddRoundConstantStage_modAdder_op2_i;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_modAdder_res_o;
  wire                SBox5Stage_SBox5Insts_0_io_input_ready;
  wire                SBox5Stage_SBox5Insts_0_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_0_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_1_io_input_ready;
  wire                SBox5Stage_SBox5Insts_1_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_1_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_2_io_input_ready;
  wire                SBox5Stage_SBox5Insts_2_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_2_io_output_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_0_payload_state_element;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_outputs_2_valid;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_2_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [4:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_7_io_inputs_0_ready;
  wire                streamMux_7_io_inputs_1_ready;
  wire                streamMux_7_io_inputs_2_ready;
  wire                streamMux_7_io_output_valid;
  wire       [6:0]    streamMux_7_io_output_payload_round_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_size;
  wire       [6:0]    streamMux_7_io_output_payload_state_id;
  wire       [254:0]  streamMux_7_io_output_payload_state_element;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_input_ready;
  wire                streamDemux_8_io_outputs_0_valid;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_0_payload_state_element;
  wire                streamDemux_8_io_outputs_1_valid;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_outputs_2_valid;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_2_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_8_io_inputs_0_ready;
  wire                streamMux_8_io_inputs_1_ready;
  wire                streamMux_8_io_inputs_2_ready;
  wire                streamMux_8_io_output_valid;
  wire       [6:0]    streamMux_8_io_output_payload_round_index;
  wire       [3:0]    streamMux_8_io_output_payload_state_size;
  wire       [6:0]    streamMux_8_io_output_payload_state_id;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_0;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_1;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_2;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_3;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_4;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_5;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_6;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_7;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_8;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_9;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_10;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_11;
  wire       [2:0]    _zz__zz_SBox5Stage_DemuxSelect_1;
  wire       [2:0]    _zz__zz_MDSMixStage_DemuxSelect_1;
  wire                AddRoundConstantStage_output_valid;
  reg                 AddRoundConstantStage_output_ready;
  wire       [6:0]    AddRoundConstantStage_output_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_payload_state_id;
  reg        [254:0]  AddRoundConstantStage_output_payload_state_element;
  wire                when_PoseidonThread_l46;
  wire                AddRoundConstantStage_output_m2sPipe_valid;
  wire                AddRoundConstantStage_output_m2sPipe_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_payload_state_element;
  reg                 AddRoundConstantStage_output_rValid;
  reg        [6:0]    AddRoundConstantStage_output_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_rData_state_element;
  wire                when_Stream_l342;
  wire                AddRoundConstantStage_output_m2sPipe_input_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_payload_state_element;
  reg                 AddRoundConstantStage_output_m2sPipe_rValid;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect_1;
  wire                _zz_SBox5Stage_DemuxSelect_2;
  wire                _zz_SBox5Stage_DemuxSelect_3;
  wire       [1:0]    SBox5Stage_DemuxSelect;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_SBox5Stage_output_valid;
  wire                _zz_io_pop_ready;
  wire                SBox5Stage_output_valid;
  reg                 SBox5Stage_output_ready;
  wire       [6:0]    SBox5Stage_output_payload_round_index;
  wire       [3:0]    SBox5Stage_output_payload_state_index;
  wire       [3:0]    SBox5Stage_output_payload_state_size;
  wire       [6:0]    SBox5Stage_output_payload_state_id;
  wire       [254:0]  SBox5Stage_output_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_valid;
  wire                SBox5Stage_output_m2sPipe_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_payload_state_element;
  reg                 SBox5Stage_output_rValid;
  reg        [6:0]    SBox5Stage_output_rData_round_index;
  reg        [3:0]    SBox5Stage_output_rData_state_index;
  reg        [3:0]    SBox5Stage_output_rData_state_size;
  reg        [6:0]    SBox5Stage_output_rData_state_id;
  reg        [254:0]  SBox5Stage_output_rData_state_element;
  wire                when_Stream_l342_1;
  wire                SBox5Stage_output_m2sPipe_input_valid;
  wire                SBox5Stage_output_m2sPipe_input_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_payload_state_element;
  reg                 SBox5Stage_output_m2sPipe_rValid;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_round_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_size;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_state_id;
  reg        [254:0]  SBox5Stage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect_1;
  wire                _zz_MDSMixStage_DemuxSelect_2;
  wire                _zz_MDSMixStage_DemuxSelect_3;
  wire       [1:0]    MDSMixStage_DemuxSelect;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_MDSMixStage_output_valid;
  wire                _zz_io_pop_ready_1;
  wire                MDSMixStage_output_valid;
  wire                MDSMixStage_output_ready;
  wire       [6:0]    MDSMixStage_output_payload_round_index;
  wire       [3:0]    MDSMixStage_output_payload_state_size;
  wire       [6:0]    MDSMixStage_output_payload_state_id;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_11;

  assign _zz__zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect - 3'b001);
  assign _zz__zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect - 3'b001);
  RoundConstants_8 AddRoundConstantStage_roundConstants_t3 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_9 AddRoundConstantStage_roundConstants_t5 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_10 AddRoundConstantStage_roundConstants_t9 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                  ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                  )  //i
  );
  RoundConstants_11 AddRoundConstantStage_roundConstants_t12 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                   ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                   )  //i
  );
  ModAdder AddRoundConstantStage_modAdder (
    .op1_i    (io_input_payload_state_element        ), //i
    .op2_i    (AddRoundConstantStage_modAdder_op2_i  ), //i
    .res_o    (AddRoundConstantStage_modAdder_res_o  )  //o
  );
  SBox5 SBox5Stage_SBox5Insts_0 (
    .io_input_valid                     (streamDemux_7_io_outputs_0_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_0_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_0_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_0_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_0_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_0_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_0_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_0_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_1 (
    .io_input_valid                     (streamDemux_7_io_outputs_1_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_1_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_1_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_1_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_1_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_1_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_1_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_1_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_2 (
    .io_input_valid                     (streamDemux_7_io_outputs_2_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_2_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_2_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_2_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_2_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_2_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_2_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_2_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  StreamFork_10 AddRoundConstantStage_output_m2sPipe_input_fork (
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_7_io_input_ready                                                        ), //i
    .io_outputs_0_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_7 (
    .io_select                             (SBox5Stage_DemuxSelect                                                              ), //i
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_7_io_input_ready                                                        ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_7_io_outputs_0_valid                                                    ), //o
    .io_outputs_0_ready                    (SBox5Stage_SBox5Insts_0_io_input_ready                                              ), //i
    .io_outputs_0_payload_round_index      (streamDemux_7_io_outputs_0_payload_round_index                                      ), //o
    .io_outputs_0_payload_state_index      (streamDemux_7_io_outputs_0_payload_state_index                                      ), //o
    .io_outputs_0_payload_state_size       (streamDemux_7_io_outputs_0_payload_state_size                                       ), //o
    .io_outputs_0_payload_state_id         (streamDemux_7_io_outputs_0_payload_state_id                                         ), //o
    .io_outputs_0_payload_state_element    (streamDemux_7_io_outputs_0_payload_state_element                                    ), //o
    .io_outputs_1_valid                    (streamDemux_7_io_outputs_1_valid                                                    ), //o
    .io_outputs_1_ready                    (SBox5Stage_SBox5Insts_1_io_input_ready                                              ), //i
    .io_outputs_1_payload_round_index      (streamDemux_7_io_outputs_1_payload_round_index                                      ), //o
    .io_outputs_1_payload_state_index      (streamDemux_7_io_outputs_1_payload_state_index                                      ), //o
    .io_outputs_1_payload_state_size       (streamDemux_7_io_outputs_1_payload_state_size                                       ), //o
    .io_outputs_1_payload_state_id         (streamDemux_7_io_outputs_1_payload_state_id                                         ), //o
    .io_outputs_1_payload_state_element    (streamDemux_7_io_outputs_1_payload_state_element                                    ), //o
    .io_outputs_2_valid                    (streamDemux_7_io_outputs_2_valid                                                    ), //o
    .io_outputs_2_ready                    (SBox5Stage_SBox5Insts_2_io_input_ready                                              ), //i
    .io_outputs_2_payload_round_index      (streamDemux_7_io_outputs_2_payload_round_index                                      ), //o
    .io_outputs_2_payload_state_index      (streamDemux_7_io_outputs_2_payload_state_index                                      ), //o
    .io_outputs_2_payload_state_size       (streamDemux_7_io_outputs_2_payload_state_size                                       ), //o
    .io_outputs_2_payload_state_id         (streamDemux_7_io_outputs_2_payload_state_id                                         ), //o
    .io_outputs_2_payload_state_element    (streamDemux_7_io_outputs_2_payload_state_element                                    )  //o
  );
  StreamFifoLowLatency AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready                                                                             ), //i
    .io_pop_payload     (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                                         ), //i
    .io_occupancy       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                                          ), //i
    .reset              (reset                                                                                        )  //i
  );
  StreamMux streamMux_7 (
    .io_select                            (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                                                      ), //i
    .io_inputs_0_ready                    (streamMux_7_io_inputs_0_ready                                                                ), //o
    .io_inputs_0_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index                                        ), //i
    .io_inputs_0_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index                                        ), //i
    .io_inputs_0_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size                                         ), //i
    .io_inputs_0_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id                                           ), //i
    .io_inputs_0_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element                                      ), //i
    .io_inputs_1_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                                                      ), //i
    .io_inputs_1_ready                    (streamMux_7_io_inputs_1_ready                                                                ), //o
    .io_inputs_1_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index                                        ), //i
    .io_inputs_1_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index                                        ), //i
    .io_inputs_1_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size                                         ), //i
    .io_inputs_1_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id                                           ), //i
    .io_inputs_1_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element                                      ), //i
    .io_inputs_2_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                                                      ), //i
    .io_inputs_2_ready                    (streamMux_7_io_inputs_2_ready                                                                ), //o
    .io_inputs_2_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index                                        ), //i
    .io_inputs_2_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index                                        ), //i
    .io_inputs_2_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size                                         ), //i
    .io_inputs_2_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id                                           ), //i
    .io_inputs_2_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element                                      ), //i
    .io_output_valid                      (streamMux_7_io_output_valid                                                                  ), //o
    .io_output_ready                      (_zz_io_pop_ready                                                                             ), //i
    .io_output_payload_round_index        (streamMux_7_io_output_payload_round_index                                                    ), //o
    .io_output_payload_state_index        (streamMux_7_io_output_payload_state_index                                                    ), //o
    .io_output_payload_state_size         (streamMux_7_io_output_payload_state_size                                                     ), //o
    .io_output_payload_state_id           (streamMux_7_io_output_payload_state_id                                                       ), //o
    .io_output_payload_state_element      (streamMux_7_io_output_payload_state_element                                                  )  //o
  );
  MDSMatrixMultiplier_6 MDSMixStage_matrixMultiplierInsts_0 (
    .io_input_valid                         (streamDemux_8_io_outputs_0_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_0_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_0_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_0_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_0_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_0_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_0_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_7 MDSMixStage_matrixMultiplierInsts_1 (
    .io_input_valid                         (streamDemux_8_io_outputs_1_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_1_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_1_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_1_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_1_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_1_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_1_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_8 MDSMixStage_matrixMultiplierInsts_2 (
    .io_input_valid                         (streamDemux_8_io_outputs_2_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_2_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_2_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_2_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_2_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_2_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_2_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  StreamFork_10 SBox5Stage_output_m2sPipe_input_fork (
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (SBox5Stage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_8_io_input_ready                                             ), //i
    .io_outputs_0_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_8 (
    .io_select                             (MDSMixStage_DemuxSelect                                                  ), //i
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_8_io_input_ready                                             ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_8_io_outputs_0_valid                                         ), //o
    .io_outputs_0_ready                    (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //i
    .io_outputs_0_payload_round_index      (streamDemux_8_io_outputs_0_payload_round_index                           ), //o
    .io_outputs_0_payload_state_index      (streamDemux_8_io_outputs_0_payload_state_index                           ), //o
    .io_outputs_0_payload_state_size       (streamDemux_8_io_outputs_0_payload_state_size                            ), //o
    .io_outputs_0_payload_state_id         (streamDemux_8_io_outputs_0_payload_state_id                              ), //o
    .io_outputs_0_payload_state_element    (streamDemux_8_io_outputs_0_payload_state_element                         ), //o
    .io_outputs_1_valid                    (streamDemux_8_io_outputs_1_valid                                         ), //o
    .io_outputs_1_ready                    (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //i
    .io_outputs_1_payload_round_index      (streamDemux_8_io_outputs_1_payload_round_index                           ), //o
    .io_outputs_1_payload_state_index      (streamDemux_8_io_outputs_1_payload_state_index                           ), //o
    .io_outputs_1_payload_state_size       (streamDemux_8_io_outputs_1_payload_state_size                            ), //o
    .io_outputs_1_payload_state_id         (streamDemux_8_io_outputs_1_payload_state_id                              ), //o
    .io_outputs_1_payload_state_element    (streamDemux_8_io_outputs_1_payload_state_element                         ), //o
    .io_outputs_2_valid                    (streamDemux_8_io_outputs_2_valid                                         ), //o
    .io_outputs_2_ready                    (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //i
    .io_outputs_2_payload_round_index      (streamDemux_8_io_outputs_2_payload_round_index                           ), //o
    .io_outputs_2_payload_state_index      (streamDemux_8_io_outputs_2_payload_state_index                           ), //o
    .io_outputs_2_payload_state_size       (streamDemux_8_io_outputs_2_payload_state_size                            ), //o
    .io_outputs_2_payload_state_id         (streamDemux_8_io_outputs_2_payload_state_id                              ), //o
    .io_outputs_2_payload_state_element    (streamDemux_8_io_outputs_2_payload_state_element                         )  //o
  );
  StreamFifoLowLatency_1 SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready_1                                                                ), //i
    .io_pop_payload     (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                              ), //i
    .io_occupancy       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                               ), //i
    .reset              (reset                                                                             )  //i
  );
  StreamMux_1 streamMux_8 (
    .io_select                                (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                               ), //i
    .io_inputs_0_ready                        (streamMux_8_io_inputs_0_ready                                                     ), //o
    .io_inputs_0_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index                 ), //i
    .io_inputs_0_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size                  ), //i
    .io_inputs_0_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id                    ), //i
    .io_inputs_0_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0            ), //i
    .io_inputs_0_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1            ), //i
    .io_inputs_0_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2            ), //i
    .io_inputs_0_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3            ), //i
    .io_inputs_0_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4            ), //i
    .io_inputs_0_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5            ), //i
    .io_inputs_0_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6            ), //i
    .io_inputs_0_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7            ), //i
    .io_inputs_0_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8            ), //i
    .io_inputs_0_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9            ), //i
    .io_inputs_0_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10           ), //i
    .io_inputs_0_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11           ), //i
    .io_inputs_1_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                               ), //i
    .io_inputs_1_ready                        (streamMux_8_io_inputs_1_ready                                                     ), //o
    .io_inputs_1_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index                 ), //i
    .io_inputs_1_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size                  ), //i
    .io_inputs_1_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id                    ), //i
    .io_inputs_1_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0            ), //i
    .io_inputs_1_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1            ), //i
    .io_inputs_1_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2            ), //i
    .io_inputs_1_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3            ), //i
    .io_inputs_1_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4            ), //i
    .io_inputs_1_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5            ), //i
    .io_inputs_1_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6            ), //i
    .io_inputs_1_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7            ), //i
    .io_inputs_1_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8            ), //i
    .io_inputs_1_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9            ), //i
    .io_inputs_1_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10           ), //i
    .io_inputs_1_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11           ), //i
    .io_inputs_2_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                               ), //i
    .io_inputs_2_ready                        (streamMux_8_io_inputs_2_ready                                                     ), //o
    .io_inputs_2_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index                 ), //i
    .io_inputs_2_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size                  ), //i
    .io_inputs_2_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id                    ), //i
    .io_inputs_2_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0            ), //i
    .io_inputs_2_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1            ), //i
    .io_inputs_2_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2            ), //i
    .io_inputs_2_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3            ), //i
    .io_inputs_2_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4            ), //i
    .io_inputs_2_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5            ), //i
    .io_inputs_2_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6            ), //i
    .io_inputs_2_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7            ), //i
    .io_inputs_2_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8            ), //i
    .io_inputs_2_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9            ), //i
    .io_inputs_2_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10           ), //i
    .io_inputs_2_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11           ), //i
    .io_output_valid                          (streamMux_8_io_output_valid                                                       ), //o
    .io_output_ready                          (_zz_io_pop_ready_1                                                                ), //i
    .io_output_payload_round_index            (streamMux_8_io_output_payload_round_index                                         ), //o
    .io_output_payload_state_size             (streamMux_8_io_output_payload_state_size                                          ), //o
    .io_output_payload_state_id               (streamMux_8_io_output_payload_state_id                                            ), //o
    .io_output_payload_state_elements_0       (streamMux_8_io_output_payload_state_elements_0                                    ), //o
    .io_output_payload_state_elements_1       (streamMux_8_io_output_payload_state_elements_1                                    ), //o
    .io_output_payload_state_elements_2       (streamMux_8_io_output_payload_state_elements_2                                    ), //o
    .io_output_payload_state_elements_3       (streamMux_8_io_output_payload_state_elements_3                                    ), //o
    .io_output_payload_state_elements_4       (streamMux_8_io_output_payload_state_elements_4                                    ), //o
    .io_output_payload_state_elements_5       (streamMux_8_io_output_payload_state_elements_5                                    ), //o
    .io_output_payload_state_elements_6       (streamMux_8_io_output_payload_state_elements_6                                    ), //o
    .io_output_payload_state_elements_7       (streamMux_8_io_output_payload_state_elements_7                                    ), //o
    .io_output_payload_state_elements_8       (streamMux_8_io_output_payload_state_elements_8                                    ), //o
    .io_output_payload_state_elements_9       (streamMux_8_io_output_payload_state_elements_9                                    ), //o
    .io_output_payload_state_elements_10      (streamMux_8_io_output_payload_state_elements_10                                   ), //o
    .io_output_payload_state_elements_11      (streamMux_8_io_output_payload_state_elements_11                                   )  //o
  );
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index = io_input_payload_state_index[1:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index = io_input_payload_state_index[2:0];
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
      end
      4'b0101 : begin
        if(when_PoseidonThread_l46) begin
          AddRoundConstantStage_modAdder_op2_i = 255'h0;
        end else begin
          AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
        end
      end
      4'b1001 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
      end
      4'b1100 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
      end
      default : begin
        AddRoundConstantStage_modAdder_op2_i = 255'h0;
      end
    endcase
  end

  assign when_PoseidonThread_l46 = (io_input_payload_state_index == 4'b0101);
  assign AddRoundConstantStage_output_valid = io_input_valid;
  assign io_input_ready = AddRoundConstantStage_output_ready;
  assign AddRoundConstantStage_output_payload_round_index = io_input_payload_round_index;
  assign AddRoundConstantStage_output_payload_state_index = io_input_payload_state_index;
  assign AddRoundConstantStage_output_payload_state_size = io_input_payload_state_size;
  assign AddRoundConstantStage_output_payload_state_id = io_input_payload_state_id;
  always @(*) begin
    AddRoundConstantStage_output_payload_state_element = io_input_payload_state_element;
    AddRoundConstantStage_output_payload_state_element = AddRoundConstantStage_modAdder_res_o;
  end

  always @(*) begin
    AddRoundConstantStage_output_ready = AddRoundConstantStage_output_m2sPipe_ready;
    if(when_Stream_l342) begin
      AddRoundConstantStage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! AddRoundConstantStage_output_m2sPipe_valid);
  assign AddRoundConstantStage_output_m2sPipe_valid = AddRoundConstantStage_output_rValid;
  assign AddRoundConstantStage_output_m2sPipe_payload_round_index = AddRoundConstantStage_output_rData_round_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_index = AddRoundConstantStage_output_rData_state_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_size = AddRoundConstantStage_output_rData_state_size;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_id = AddRoundConstantStage_output_rData_state_id;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_element = AddRoundConstantStage_output_rData_state_element;
  assign AddRoundConstantStage_output_m2sPipe_ready = (! AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_valid = (AddRoundConstantStage_output_m2sPipe_valid || AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_round_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_round_index : AddRoundConstantStage_output_m2sPipe_payload_round_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_index : AddRoundConstantStage_output_m2sPipe_payload_state_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_size = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_size : AddRoundConstantStage_output_m2sPipe_payload_state_size);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_id = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_id : AddRoundConstantStage_output_m2sPipe_payload_state_id);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_element = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_element : AddRoundConstantStage_output_m2sPipe_payload_state_element);
  assign AddRoundConstantStage_output_m2sPipe_input_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_SBox5Stage_DemuxSelect = {SBox5Stage_SBox5Insts_2_io_input_ready,{SBox5Stage_SBox5Insts_1_io_input_ready,SBox5Stage_SBox5Insts_0_io_input_ready}};
  assign _zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect & (~ _zz__zz_SBox5Stage_DemuxSelect_1));
  assign _zz_SBox5Stage_DemuxSelect_2 = _zz_SBox5Stage_DemuxSelect_1[1];
  assign _zz_SBox5Stage_DemuxSelect_3 = _zz_SBox5Stage_DemuxSelect_1[2];
  assign SBox5Stage_DemuxSelect = {_zz_SBox5Stage_DemuxSelect_3,_zz_SBox5Stage_DemuxSelect_2};
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = SBox5Stage_DemuxSelect;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready = (_zz_SBox5Stage_output_valid && SBox5Stage_output_ready);
  assign _zz_SBox5Stage_output_valid = (streamMux_7_io_output_valid && AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign SBox5Stage_output_valid = _zz_SBox5Stage_output_valid;
  assign SBox5Stage_output_payload_round_index = streamMux_7_io_output_payload_round_index;
  assign SBox5Stage_output_payload_state_index = streamMux_7_io_output_payload_state_index;
  assign SBox5Stage_output_payload_state_size = streamMux_7_io_output_payload_state_size;
  assign SBox5Stage_output_payload_state_id = streamMux_7_io_output_payload_state_id;
  assign SBox5Stage_output_payload_state_element = streamMux_7_io_output_payload_state_element;
  always @(*) begin
    SBox5Stage_output_ready = SBox5Stage_output_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      SBox5Stage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! SBox5Stage_output_m2sPipe_valid);
  assign SBox5Stage_output_m2sPipe_valid = SBox5Stage_output_rValid;
  assign SBox5Stage_output_m2sPipe_payload_round_index = SBox5Stage_output_rData_round_index;
  assign SBox5Stage_output_m2sPipe_payload_state_index = SBox5Stage_output_rData_state_index;
  assign SBox5Stage_output_m2sPipe_payload_state_size = SBox5Stage_output_rData_state_size;
  assign SBox5Stage_output_m2sPipe_payload_state_id = SBox5Stage_output_rData_state_id;
  assign SBox5Stage_output_m2sPipe_payload_state_element = SBox5Stage_output_rData_state_element;
  assign SBox5Stage_output_m2sPipe_ready = (! SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_valid = (SBox5Stage_output_m2sPipe_valid || SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_payload_round_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_round_index : SBox5Stage_output_m2sPipe_payload_round_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_index : SBox5Stage_output_m2sPipe_payload_state_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_size = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_size : SBox5Stage_output_m2sPipe_payload_state_size);
  assign SBox5Stage_output_m2sPipe_input_payload_state_id = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_id : SBox5Stage_output_m2sPipe_payload_state_id);
  assign SBox5Stage_output_m2sPipe_input_payload_state_element = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_element : SBox5Stage_output_m2sPipe_payload_state_element);
  assign SBox5Stage_output_m2sPipe_input_ready = SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_MDSMixStage_DemuxSelect = {MDSMixStage_matrixMultiplierInsts_2_io_input_ready,{MDSMixStage_matrixMultiplierInsts_1_io_input_ready,MDSMixStage_matrixMultiplierInsts_0_io_input_ready}};
  assign _zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect & (~ _zz__zz_MDSMixStage_DemuxSelect_1));
  assign _zz_MDSMixStage_DemuxSelect_2 = _zz_MDSMixStage_DemuxSelect_1[1];
  assign _zz_MDSMixStage_DemuxSelect_3 = _zz_MDSMixStage_DemuxSelect_1[2];
  assign MDSMixStage_DemuxSelect = {_zz_MDSMixStage_DemuxSelect_3,_zz_MDSMixStage_DemuxSelect_2};
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = MDSMixStage_DemuxSelect;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready_1 = (_zz_MDSMixStage_output_valid && MDSMixStage_output_ready);
  assign _zz_MDSMixStage_output_valid = (streamMux_8_io_output_valid && SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign MDSMixStage_output_valid = _zz_MDSMixStage_output_valid;
  assign MDSMixStage_output_payload_round_index = streamMux_8_io_output_payload_round_index;
  assign MDSMixStage_output_payload_state_size = streamMux_8_io_output_payload_state_size;
  assign MDSMixStage_output_payload_state_id = streamMux_8_io_output_payload_state_id;
  assign MDSMixStage_output_payload_state_elements_0 = streamMux_8_io_output_payload_state_elements_0;
  assign MDSMixStage_output_payload_state_elements_1 = streamMux_8_io_output_payload_state_elements_1;
  assign MDSMixStage_output_payload_state_elements_2 = streamMux_8_io_output_payload_state_elements_2;
  assign MDSMixStage_output_payload_state_elements_3 = streamMux_8_io_output_payload_state_elements_3;
  assign MDSMixStage_output_payload_state_elements_4 = streamMux_8_io_output_payload_state_elements_4;
  assign MDSMixStage_output_payload_state_elements_5 = streamMux_8_io_output_payload_state_elements_5;
  assign MDSMixStage_output_payload_state_elements_6 = streamMux_8_io_output_payload_state_elements_6;
  assign MDSMixStage_output_payload_state_elements_7 = streamMux_8_io_output_payload_state_elements_7;
  assign MDSMixStage_output_payload_state_elements_8 = streamMux_8_io_output_payload_state_elements_8;
  assign MDSMixStage_output_payload_state_elements_9 = streamMux_8_io_output_payload_state_elements_9;
  assign MDSMixStage_output_payload_state_elements_10 = streamMux_8_io_output_payload_state_elements_10;
  assign MDSMixStage_output_payload_state_elements_11 = streamMux_8_io_output_payload_state_elements_11;
  assign io_output_valid = MDSMixStage_output_valid;
  assign MDSMixStage_output_ready = io_output_ready;
  assign io_output_payload_round_index = MDSMixStage_output_payload_round_index;
  assign io_output_payload_state_size = MDSMixStage_output_payload_state_size;
  assign io_output_payload_state_id = MDSMixStage_output_payload_state_id;
  assign io_output_payload_state_elements_0 = MDSMixStage_output_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = MDSMixStage_output_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = MDSMixStage_output_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = MDSMixStage_output_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = MDSMixStage_output_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = MDSMixStage_output_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = MDSMixStage_output_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = MDSMixStage_output_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = MDSMixStage_output_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = MDSMixStage_output_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = MDSMixStage_output_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = MDSMixStage_output_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      AddRoundConstantStage_output_rValid <= 1'b0;
      AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      SBox5Stage_output_rValid <= 1'b0;
      SBox5Stage_output_m2sPipe_rValid <= 1'b0;
    end else begin
      if(AddRoundConstantStage_output_ready) begin
        AddRoundConstantStage_output_rValid <= AddRoundConstantStage_output_valid;
      end
      if(AddRoundConstantStage_output_m2sPipe_valid) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b1;
      end
      if(AddRoundConstantStage_output_m2sPipe_input_ready) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      end
      if(SBox5Stage_output_ready) begin
        SBox5Stage_output_rValid <= SBox5Stage_output_valid;
      end
      if(SBox5Stage_output_m2sPipe_valid) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b1;
      end
      if(SBox5Stage_output_m2sPipe_input_ready) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(AddRoundConstantStage_output_ready) begin
      AddRoundConstantStage_output_rData_round_index <= AddRoundConstantStage_output_payload_round_index;
      AddRoundConstantStage_output_rData_state_index <= AddRoundConstantStage_output_payload_state_index;
      AddRoundConstantStage_output_rData_state_size <= AddRoundConstantStage_output_payload_state_size;
      AddRoundConstantStage_output_rData_state_id <= AddRoundConstantStage_output_payload_state_id;
      AddRoundConstantStage_output_rData_state_element <= AddRoundConstantStage_output_payload_state_element;
    end
    if(AddRoundConstantStage_output_m2sPipe_ready) begin
      AddRoundConstantStage_output_m2sPipe_rData_round_index <= AddRoundConstantStage_output_m2sPipe_payload_round_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_index <= AddRoundConstantStage_output_m2sPipe_payload_state_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_size <= AddRoundConstantStage_output_m2sPipe_payload_state_size;
      AddRoundConstantStage_output_m2sPipe_rData_state_id <= AddRoundConstantStage_output_m2sPipe_payload_state_id;
      AddRoundConstantStage_output_m2sPipe_rData_state_element <= AddRoundConstantStage_output_m2sPipe_payload_state_element;
    end
    if(SBox5Stage_output_ready) begin
      SBox5Stage_output_rData_round_index <= SBox5Stage_output_payload_round_index;
      SBox5Stage_output_rData_state_index <= SBox5Stage_output_payload_state_index;
      SBox5Stage_output_rData_state_size <= SBox5Stage_output_payload_state_size;
      SBox5Stage_output_rData_state_id <= SBox5Stage_output_payload_state_id;
      SBox5Stage_output_rData_state_element <= SBox5Stage_output_payload_state_element;
    end
    if(SBox5Stage_output_m2sPipe_ready) begin
      SBox5Stage_output_m2sPipe_rData_round_index <= SBox5Stage_output_m2sPipe_payload_round_index;
      SBox5Stage_output_m2sPipe_rData_state_index <= SBox5Stage_output_m2sPipe_payload_state_index;
      SBox5Stage_output_m2sPipe_rData_state_size <= SBox5Stage_output_m2sPipe_payload_state_size;
      SBox5Stage_output_m2sPipe_rData_state_id <= SBox5Stage_output_m2sPipe_payload_state_id;
      SBox5Stage_output_m2sPipe_rData_state_element <= SBox5Stage_output_m2sPipe_payload_state_element;
    end
  end


endmodule

module PoseidonThread_1 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index;
  wire       [2:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index;
  reg        [254:0]  AddRoundConstantStage_modAdder_op2_i;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_modAdder_res_o;
  wire                SBox5Stage_SBox5Insts_0_io_input_ready;
  wire                SBox5Stage_SBox5Insts_0_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_0_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_1_io_input_ready;
  wire                SBox5Stage_SBox5Insts_1_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_1_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_2_io_input_ready;
  wire                SBox5Stage_SBox5Insts_2_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_2_io_output_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_0_payload_state_element;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_outputs_2_valid;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_2_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [4:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_7_io_inputs_0_ready;
  wire                streamMux_7_io_inputs_1_ready;
  wire                streamMux_7_io_inputs_2_ready;
  wire                streamMux_7_io_output_valid;
  wire       [6:0]    streamMux_7_io_output_payload_round_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_size;
  wire       [6:0]    streamMux_7_io_output_payload_state_id;
  wire       [254:0]  streamMux_7_io_output_payload_state_element;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_input_ready;
  wire                streamDemux_8_io_outputs_0_valid;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_0_payload_state_element;
  wire                streamDemux_8_io_outputs_1_valid;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_outputs_2_valid;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_2_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_8_io_inputs_0_ready;
  wire                streamMux_8_io_inputs_1_ready;
  wire                streamMux_8_io_inputs_2_ready;
  wire                streamMux_8_io_output_valid;
  wire       [6:0]    streamMux_8_io_output_payload_round_index;
  wire       [3:0]    streamMux_8_io_output_payload_state_size;
  wire       [6:0]    streamMux_8_io_output_payload_state_id;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_0;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_1;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_2;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_3;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_4;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_5;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_6;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_7;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_8;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_9;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_10;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_11;
  wire       [2:0]    _zz__zz_SBox5Stage_DemuxSelect_1;
  wire       [2:0]    _zz__zz_MDSMixStage_DemuxSelect_1;
  wire                AddRoundConstantStage_output_valid;
  reg                 AddRoundConstantStage_output_ready;
  wire       [6:0]    AddRoundConstantStage_output_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_payload_state_id;
  reg        [254:0]  AddRoundConstantStage_output_payload_state_element;
  wire                when_PoseidonThread_l46;
  wire                AddRoundConstantStage_output_m2sPipe_valid;
  wire                AddRoundConstantStage_output_m2sPipe_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_payload_state_element;
  reg                 AddRoundConstantStage_output_rValid;
  reg        [6:0]    AddRoundConstantStage_output_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_rData_state_element;
  wire                when_Stream_l342;
  wire                AddRoundConstantStage_output_m2sPipe_input_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_payload_state_element;
  reg                 AddRoundConstantStage_output_m2sPipe_rValid;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect_1;
  wire                _zz_SBox5Stage_DemuxSelect_2;
  wire                _zz_SBox5Stage_DemuxSelect_3;
  wire       [1:0]    SBox5Stage_DemuxSelect;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_SBox5Stage_output_valid;
  wire                _zz_io_pop_ready;
  wire                SBox5Stage_output_valid;
  reg                 SBox5Stage_output_ready;
  wire       [6:0]    SBox5Stage_output_payload_round_index;
  wire       [3:0]    SBox5Stage_output_payload_state_index;
  wire       [3:0]    SBox5Stage_output_payload_state_size;
  wire       [6:0]    SBox5Stage_output_payload_state_id;
  wire       [254:0]  SBox5Stage_output_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_valid;
  wire                SBox5Stage_output_m2sPipe_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_payload_state_element;
  reg                 SBox5Stage_output_rValid;
  reg        [6:0]    SBox5Stage_output_rData_round_index;
  reg        [3:0]    SBox5Stage_output_rData_state_index;
  reg        [3:0]    SBox5Stage_output_rData_state_size;
  reg        [6:0]    SBox5Stage_output_rData_state_id;
  reg        [254:0]  SBox5Stage_output_rData_state_element;
  wire                when_Stream_l342_1;
  wire                SBox5Stage_output_m2sPipe_input_valid;
  wire                SBox5Stage_output_m2sPipe_input_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_payload_state_element;
  reg                 SBox5Stage_output_m2sPipe_rValid;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_round_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_size;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_state_id;
  reg        [254:0]  SBox5Stage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect_1;
  wire                _zz_MDSMixStage_DemuxSelect_2;
  wire                _zz_MDSMixStage_DemuxSelect_3;
  wire       [1:0]    MDSMixStage_DemuxSelect;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_MDSMixStage_output_valid;
  wire                _zz_io_pop_ready_1;
  wire                MDSMixStage_output_valid;
  wire                MDSMixStage_output_ready;
  wire       [6:0]    MDSMixStage_output_payload_round_index;
  wire       [3:0]    MDSMixStage_output_payload_state_size;
  wire       [6:0]    MDSMixStage_output_payload_state_id;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_11;

  assign _zz__zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect - 3'b001);
  assign _zz__zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect - 3'b001);
  RoundConstants_4 AddRoundConstantStage_roundConstants_t3 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_5 AddRoundConstantStage_roundConstants_t5 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_6 AddRoundConstantStage_roundConstants_t9 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                  ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                  )  //i
  );
  RoundConstants_7 AddRoundConstantStage_roundConstants_t12 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                   ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                   )  //i
  );
  ModAdder AddRoundConstantStage_modAdder (
    .op1_i    (io_input_payload_state_element        ), //i
    .op2_i    (AddRoundConstantStage_modAdder_op2_i  ), //i
    .res_o    (AddRoundConstantStage_modAdder_res_o  )  //o
  );
  SBox5 SBox5Stage_SBox5Insts_0 (
    .io_input_valid                     (streamDemux_7_io_outputs_0_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_0_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_0_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_0_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_0_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_0_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_0_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_0_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_1 (
    .io_input_valid                     (streamDemux_7_io_outputs_1_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_1_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_1_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_1_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_1_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_1_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_1_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_1_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_2 (
    .io_input_valid                     (streamDemux_7_io_outputs_2_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_2_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_2_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_2_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_2_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_2_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_2_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_2_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  StreamFork_10 AddRoundConstantStage_output_m2sPipe_input_fork (
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_7_io_input_ready                                                        ), //i
    .io_outputs_0_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_7 (
    .io_select                             (SBox5Stage_DemuxSelect                                                              ), //i
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_7_io_input_ready                                                        ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_7_io_outputs_0_valid                                                    ), //o
    .io_outputs_0_ready                    (SBox5Stage_SBox5Insts_0_io_input_ready                                              ), //i
    .io_outputs_0_payload_round_index      (streamDemux_7_io_outputs_0_payload_round_index                                      ), //o
    .io_outputs_0_payload_state_index      (streamDemux_7_io_outputs_0_payload_state_index                                      ), //o
    .io_outputs_0_payload_state_size       (streamDemux_7_io_outputs_0_payload_state_size                                       ), //o
    .io_outputs_0_payload_state_id         (streamDemux_7_io_outputs_0_payload_state_id                                         ), //o
    .io_outputs_0_payload_state_element    (streamDemux_7_io_outputs_0_payload_state_element                                    ), //o
    .io_outputs_1_valid                    (streamDemux_7_io_outputs_1_valid                                                    ), //o
    .io_outputs_1_ready                    (SBox5Stage_SBox5Insts_1_io_input_ready                                              ), //i
    .io_outputs_1_payload_round_index      (streamDemux_7_io_outputs_1_payload_round_index                                      ), //o
    .io_outputs_1_payload_state_index      (streamDemux_7_io_outputs_1_payload_state_index                                      ), //o
    .io_outputs_1_payload_state_size       (streamDemux_7_io_outputs_1_payload_state_size                                       ), //o
    .io_outputs_1_payload_state_id         (streamDemux_7_io_outputs_1_payload_state_id                                         ), //o
    .io_outputs_1_payload_state_element    (streamDemux_7_io_outputs_1_payload_state_element                                    ), //o
    .io_outputs_2_valid                    (streamDemux_7_io_outputs_2_valid                                                    ), //o
    .io_outputs_2_ready                    (SBox5Stage_SBox5Insts_2_io_input_ready                                              ), //i
    .io_outputs_2_payload_round_index      (streamDemux_7_io_outputs_2_payload_round_index                                      ), //o
    .io_outputs_2_payload_state_index      (streamDemux_7_io_outputs_2_payload_state_index                                      ), //o
    .io_outputs_2_payload_state_size       (streamDemux_7_io_outputs_2_payload_state_size                                       ), //o
    .io_outputs_2_payload_state_id         (streamDemux_7_io_outputs_2_payload_state_id                                         ), //o
    .io_outputs_2_payload_state_element    (streamDemux_7_io_outputs_2_payload_state_element                                    )  //o
  );
  StreamFifoLowLatency AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready                                                                             ), //i
    .io_pop_payload     (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                                         ), //i
    .io_occupancy       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                                          ), //i
    .reset              (reset                                                                                        )  //i
  );
  StreamMux streamMux_7 (
    .io_select                            (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                                                      ), //i
    .io_inputs_0_ready                    (streamMux_7_io_inputs_0_ready                                                                ), //o
    .io_inputs_0_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index                                        ), //i
    .io_inputs_0_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index                                        ), //i
    .io_inputs_0_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size                                         ), //i
    .io_inputs_0_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id                                           ), //i
    .io_inputs_0_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element                                      ), //i
    .io_inputs_1_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                                                      ), //i
    .io_inputs_1_ready                    (streamMux_7_io_inputs_1_ready                                                                ), //o
    .io_inputs_1_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index                                        ), //i
    .io_inputs_1_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index                                        ), //i
    .io_inputs_1_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size                                         ), //i
    .io_inputs_1_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id                                           ), //i
    .io_inputs_1_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element                                      ), //i
    .io_inputs_2_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                                                      ), //i
    .io_inputs_2_ready                    (streamMux_7_io_inputs_2_ready                                                                ), //o
    .io_inputs_2_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index                                        ), //i
    .io_inputs_2_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index                                        ), //i
    .io_inputs_2_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size                                         ), //i
    .io_inputs_2_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id                                           ), //i
    .io_inputs_2_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element                                      ), //i
    .io_output_valid                      (streamMux_7_io_output_valid                                                                  ), //o
    .io_output_ready                      (_zz_io_pop_ready                                                                             ), //i
    .io_output_payload_round_index        (streamMux_7_io_output_payload_round_index                                                    ), //o
    .io_output_payload_state_index        (streamMux_7_io_output_payload_state_index                                                    ), //o
    .io_output_payload_state_size         (streamMux_7_io_output_payload_state_size                                                     ), //o
    .io_output_payload_state_id           (streamMux_7_io_output_payload_state_id                                                       ), //o
    .io_output_payload_state_element      (streamMux_7_io_output_payload_state_element                                                  )  //o
  );
  MDSMatrixMultiplier_3 MDSMixStage_matrixMultiplierInsts_0 (
    .io_input_valid                         (streamDemux_8_io_outputs_0_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_0_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_0_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_0_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_0_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_0_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_0_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_4 MDSMixStage_matrixMultiplierInsts_1 (
    .io_input_valid                         (streamDemux_8_io_outputs_1_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_1_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_1_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_1_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_1_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_1_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_1_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_5 MDSMixStage_matrixMultiplierInsts_2 (
    .io_input_valid                         (streamDemux_8_io_outputs_2_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_2_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_2_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_2_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_2_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_2_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_2_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  StreamFork_10 SBox5Stage_output_m2sPipe_input_fork (
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (SBox5Stage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_8_io_input_ready                                             ), //i
    .io_outputs_0_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_8 (
    .io_select                             (MDSMixStage_DemuxSelect                                                  ), //i
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_8_io_input_ready                                             ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_8_io_outputs_0_valid                                         ), //o
    .io_outputs_0_ready                    (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //i
    .io_outputs_0_payload_round_index      (streamDemux_8_io_outputs_0_payload_round_index                           ), //o
    .io_outputs_0_payload_state_index      (streamDemux_8_io_outputs_0_payload_state_index                           ), //o
    .io_outputs_0_payload_state_size       (streamDemux_8_io_outputs_0_payload_state_size                            ), //o
    .io_outputs_0_payload_state_id         (streamDemux_8_io_outputs_0_payload_state_id                              ), //o
    .io_outputs_0_payload_state_element    (streamDemux_8_io_outputs_0_payload_state_element                         ), //o
    .io_outputs_1_valid                    (streamDemux_8_io_outputs_1_valid                                         ), //o
    .io_outputs_1_ready                    (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //i
    .io_outputs_1_payload_round_index      (streamDemux_8_io_outputs_1_payload_round_index                           ), //o
    .io_outputs_1_payload_state_index      (streamDemux_8_io_outputs_1_payload_state_index                           ), //o
    .io_outputs_1_payload_state_size       (streamDemux_8_io_outputs_1_payload_state_size                            ), //o
    .io_outputs_1_payload_state_id         (streamDemux_8_io_outputs_1_payload_state_id                              ), //o
    .io_outputs_1_payload_state_element    (streamDemux_8_io_outputs_1_payload_state_element                         ), //o
    .io_outputs_2_valid                    (streamDemux_8_io_outputs_2_valid                                         ), //o
    .io_outputs_2_ready                    (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //i
    .io_outputs_2_payload_round_index      (streamDemux_8_io_outputs_2_payload_round_index                           ), //o
    .io_outputs_2_payload_state_index      (streamDemux_8_io_outputs_2_payload_state_index                           ), //o
    .io_outputs_2_payload_state_size       (streamDemux_8_io_outputs_2_payload_state_size                            ), //o
    .io_outputs_2_payload_state_id         (streamDemux_8_io_outputs_2_payload_state_id                              ), //o
    .io_outputs_2_payload_state_element    (streamDemux_8_io_outputs_2_payload_state_element                         )  //o
  );
  StreamFifoLowLatency_1 SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready_1                                                                ), //i
    .io_pop_payload     (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                              ), //i
    .io_occupancy       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                               ), //i
    .reset              (reset                                                                             )  //i
  );
  StreamMux_1 streamMux_8 (
    .io_select                                (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                               ), //i
    .io_inputs_0_ready                        (streamMux_8_io_inputs_0_ready                                                     ), //o
    .io_inputs_0_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index                 ), //i
    .io_inputs_0_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size                  ), //i
    .io_inputs_0_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id                    ), //i
    .io_inputs_0_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0            ), //i
    .io_inputs_0_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1            ), //i
    .io_inputs_0_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2            ), //i
    .io_inputs_0_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3            ), //i
    .io_inputs_0_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4            ), //i
    .io_inputs_0_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5            ), //i
    .io_inputs_0_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6            ), //i
    .io_inputs_0_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7            ), //i
    .io_inputs_0_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8            ), //i
    .io_inputs_0_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9            ), //i
    .io_inputs_0_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10           ), //i
    .io_inputs_0_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11           ), //i
    .io_inputs_1_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                               ), //i
    .io_inputs_1_ready                        (streamMux_8_io_inputs_1_ready                                                     ), //o
    .io_inputs_1_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index                 ), //i
    .io_inputs_1_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size                  ), //i
    .io_inputs_1_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id                    ), //i
    .io_inputs_1_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0            ), //i
    .io_inputs_1_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1            ), //i
    .io_inputs_1_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2            ), //i
    .io_inputs_1_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3            ), //i
    .io_inputs_1_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4            ), //i
    .io_inputs_1_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5            ), //i
    .io_inputs_1_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6            ), //i
    .io_inputs_1_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7            ), //i
    .io_inputs_1_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8            ), //i
    .io_inputs_1_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9            ), //i
    .io_inputs_1_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10           ), //i
    .io_inputs_1_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11           ), //i
    .io_inputs_2_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                               ), //i
    .io_inputs_2_ready                        (streamMux_8_io_inputs_2_ready                                                     ), //o
    .io_inputs_2_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index                 ), //i
    .io_inputs_2_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size                  ), //i
    .io_inputs_2_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id                    ), //i
    .io_inputs_2_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0            ), //i
    .io_inputs_2_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1            ), //i
    .io_inputs_2_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2            ), //i
    .io_inputs_2_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3            ), //i
    .io_inputs_2_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4            ), //i
    .io_inputs_2_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5            ), //i
    .io_inputs_2_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6            ), //i
    .io_inputs_2_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7            ), //i
    .io_inputs_2_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8            ), //i
    .io_inputs_2_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9            ), //i
    .io_inputs_2_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10           ), //i
    .io_inputs_2_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11           ), //i
    .io_output_valid                          (streamMux_8_io_output_valid                                                       ), //o
    .io_output_ready                          (_zz_io_pop_ready_1                                                                ), //i
    .io_output_payload_round_index            (streamMux_8_io_output_payload_round_index                                         ), //o
    .io_output_payload_state_size             (streamMux_8_io_output_payload_state_size                                          ), //o
    .io_output_payload_state_id               (streamMux_8_io_output_payload_state_id                                            ), //o
    .io_output_payload_state_elements_0       (streamMux_8_io_output_payload_state_elements_0                                    ), //o
    .io_output_payload_state_elements_1       (streamMux_8_io_output_payload_state_elements_1                                    ), //o
    .io_output_payload_state_elements_2       (streamMux_8_io_output_payload_state_elements_2                                    ), //o
    .io_output_payload_state_elements_3       (streamMux_8_io_output_payload_state_elements_3                                    ), //o
    .io_output_payload_state_elements_4       (streamMux_8_io_output_payload_state_elements_4                                    ), //o
    .io_output_payload_state_elements_5       (streamMux_8_io_output_payload_state_elements_5                                    ), //o
    .io_output_payload_state_elements_6       (streamMux_8_io_output_payload_state_elements_6                                    ), //o
    .io_output_payload_state_elements_7       (streamMux_8_io_output_payload_state_elements_7                                    ), //o
    .io_output_payload_state_elements_8       (streamMux_8_io_output_payload_state_elements_8                                    ), //o
    .io_output_payload_state_elements_9       (streamMux_8_io_output_payload_state_elements_9                                    ), //o
    .io_output_payload_state_elements_10      (streamMux_8_io_output_payload_state_elements_10                                   ), //o
    .io_output_payload_state_elements_11      (streamMux_8_io_output_payload_state_elements_11                                   )  //o
  );
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index = io_input_payload_state_index[1:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index = io_input_payload_state_index[2:0];
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
      end
      4'b0101 : begin
        if(when_PoseidonThread_l46) begin
          AddRoundConstantStage_modAdder_op2_i = 255'h0;
        end else begin
          AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
        end
      end
      4'b1001 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
      end
      4'b1100 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
      end
      default : begin
        AddRoundConstantStage_modAdder_op2_i = 255'h0;
      end
    endcase
  end

  assign when_PoseidonThread_l46 = (io_input_payload_state_index == 4'b0101);
  assign AddRoundConstantStage_output_valid = io_input_valid;
  assign io_input_ready = AddRoundConstantStage_output_ready;
  assign AddRoundConstantStage_output_payload_round_index = io_input_payload_round_index;
  assign AddRoundConstantStage_output_payload_state_index = io_input_payload_state_index;
  assign AddRoundConstantStage_output_payload_state_size = io_input_payload_state_size;
  assign AddRoundConstantStage_output_payload_state_id = io_input_payload_state_id;
  always @(*) begin
    AddRoundConstantStage_output_payload_state_element = io_input_payload_state_element;
    AddRoundConstantStage_output_payload_state_element = AddRoundConstantStage_modAdder_res_o;
  end

  always @(*) begin
    AddRoundConstantStage_output_ready = AddRoundConstantStage_output_m2sPipe_ready;
    if(when_Stream_l342) begin
      AddRoundConstantStage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! AddRoundConstantStage_output_m2sPipe_valid);
  assign AddRoundConstantStage_output_m2sPipe_valid = AddRoundConstantStage_output_rValid;
  assign AddRoundConstantStage_output_m2sPipe_payload_round_index = AddRoundConstantStage_output_rData_round_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_index = AddRoundConstantStage_output_rData_state_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_size = AddRoundConstantStage_output_rData_state_size;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_id = AddRoundConstantStage_output_rData_state_id;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_element = AddRoundConstantStage_output_rData_state_element;
  assign AddRoundConstantStage_output_m2sPipe_ready = (! AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_valid = (AddRoundConstantStage_output_m2sPipe_valid || AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_round_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_round_index : AddRoundConstantStage_output_m2sPipe_payload_round_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_index : AddRoundConstantStage_output_m2sPipe_payload_state_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_size = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_size : AddRoundConstantStage_output_m2sPipe_payload_state_size);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_id = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_id : AddRoundConstantStage_output_m2sPipe_payload_state_id);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_element = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_element : AddRoundConstantStage_output_m2sPipe_payload_state_element);
  assign AddRoundConstantStage_output_m2sPipe_input_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_SBox5Stage_DemuxSelect = {SBox5Stage_SBox5Insts_2_io_input_ready,{SBox5Stage_SBox5Insts_1_io_input_ready,SBox5Stage_SBox5Insts_0_io_input_ready}};
  assign _zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect & (~ _zz__zz_SBox5Stage_DemuxSelect_1));
  assign _zz_SBox5Stage_DemuxSelect_2 = _zz_SBox5Stage_DemuxSelect_1[1];
  assign _zz_SBox5Stage_DemuxSelect_3 = _zz_SBox5Stage_DemuxSelect_1[2];
  assign SBox5Stage_DemuxSelect = {_zz_SBox5Stage_DemuxSelect_3,_zz_SBox5Stage_DemuxSelect_2};
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = SBox5Stage_DemuxSelect;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready = (_zz_SBox5Stage_output_valid && SBox5Stage_output_ready);
  assign _zz_SBox5Stage_output_valid = (streamMux_7_io_output_valid && AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign SBox5Stage_output_valid = _zz_SBox5Stage_output_valid;
  assign SBox5Stage_output_payload_round_index = streamMux_7_io_output_payload_round_index;
  assign SBox5Stage_output_payload_state_index = streamMux_7_io_output_payload_state_index;
  assign SBox5Stage_output_payload_state_size = streamMux_7_io_output_payload_state_size;
  assign SBox5Stage_output_payload_state_id = streamMux_7_io_output_payload_state_id;
  assign SBox5Stage_output_payload_state_element = streamMux_7_io_output_payload_state_element;
  always @(*) begin
    SBox5Stage_output_ready = SBox5Stage_output_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      SBox5Stage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! SBox5Stage_output_m2sPipe_valid);
  assign SBox5Stage_output_m2sPipe_valid = SBox5Stage_output_rValid;
  assign SBox5Stage_output_m2sPipe_payload_round_index = SBox5Stage_output_rData_round_index;
  assign SBox5Stage_output_m2sPipe_payload_state_index = SBox5Stage_output_rData_state_index;
  assign SBox5Stage_output_m2sPipe_payload_state_size = SBox5Stage_output_rData_state_size;
  assign SBox5Stage_output_m2sPipe_payload_state_id = SBox5Stage_output_rData_state_id;
  assign SBox5Stage_output_m2sPipe_payload_state_element = SBox5Stage_output_rData_state_element;
  assign SBox5Stage_output_m2sPipe_ready = (! SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_valid = (SBox5Stage_output_m2sPipe_valid || SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_payload_round_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_round_index : SBox5Stage_output_m2sPipe_payload_round_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_index : SBox5Stage_output_m2sPipe_payload_state_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_size = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_size : SBox5Stage_output_m2sPipe_payload_state_size);
  assign SBox5Stage_output_m2sPipe_input_payload_state_id = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_id : SBox5Stage_output_m2sPipe_payload_state_id);
  assign SBox5Stage_output_m2sPipe_input_payload_state_element = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_element : SBox5Stage_output_m2sPipe_payload_state_element);
  assign SBox5Stage_output_m2sPipe_input_ready = SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_MDSMixStage_DemuxSelect = {MDSMixStage_matrixMultiplierInsts_2_io_input_ready,{MDSMixStage_matrixMultiplierInsts_1_io_input_ready,MDSMixStage_matrixMultiplierInsts_0_io_input_ready}};
  assign _zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect & (~ _zz__zz_MDSMixStage_DemuxSelect_1));
  assign _zz_MDSMixStage_DemuxSelect_2 = _zz_MDSMixStage_DemuxSelect_1[1];
  assign _zz_MDSMixStage_DemuxSelect_3 = _zz_MDSMixStage_DemuxSelect_1[2];
  assign MDSMixStage_DemuxSelect = {_zz_MDSMixStage_DemuxSelect_3,_zz_MDSMixStage_DemuxSelect_2};
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = MDSMixStage_DemuxSelect;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready_1 = (_zz_MDSMixStage_output_valid && MDSMixStage_output_ready);
  assign _zz_MDSMixStage_output_valid = (streamMux_8_io_output_valid && SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign MDSMixStage_output_valid = _zz_MDSMixStage_output_valid;
  assign MDSMixStage_output_payload_round_index = streamMux_8_io_output_payload_round_index;
  assign MDSMixStage_output_payload_state_size = streamMux_8_io_output_payload_state_size;
  assign MDSMixStage_output_payload_state_id = streamMux_8_io_output_payload_state_id;
  assign MDSMixStage_output_payload_state_elements_0 = streamMux_8_io_output_payload_state_elements_0;
  assign MDSMixStage_output_payload_state_elements_1 = streamMux_8_io_output_payload_state_elements_1;
  assign MDSMixStage_output_payload_state_elements_2 = streamMux_8_io_output_payload_state_elements_2;
  assign MDSMixStage_output_payload_state_elements_3 = streamMux_8_io_output_payload_state_elements_3;
  assign MDSMixStage_output_payload_state_elements_4 = streamMux_8_io_output_payload_state_elements_4;
  assign MDSMixStage_output_payload_state_elements_5 = streamMux_8_io_output_payload_state_elements_5;
  assign MDSMixStage_output_payload_state_elements_6 = streamMux_8_io_output_payload_state_elements_6;
  assign MDSMixStage_output_payload_state_elements_7 = streamMux_8_io_output_payload_state_elements_7;
  assign MDSMixStage_output_payload_state_elements_8 = streamMux_8_io_output_payload_state_elements_8;
  assign MDSMixStage_output_payload_state_elements_9 = streamMux_8_io_output_payload_state_elements_9;
  assign MDSMixStage_output_payload_state_elements_10 = streamMux_8_io_output_payload_state_elements_10;
  assign MDSMixStage_output_payload_state_elements_11 = streamMux_8_io_output_payload_state_elements_11;
  assign io_output_valid = MDSMixStage_output_valid;
  assign MDSMixStage_output_ready = io_output_ready;
  assign io_output_payload_round_index = MDSMixStage_output_payload_round_index;
  assign io_output_payload_state_size = MDSMixStage_output_payload_state_size;
  assign io_output_payload_state_id = MDSMixStage_output_payload_state_id;
  assign io_output_payload_state_elements_0 = MDSMixStage_output_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = MDSMixStage_output_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = MDSMixStage_output_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = MDSMixStage_output_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = MDSMixStage_output_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = MDSMixStage_output_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = MDSMixStage_output_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = MDSMixStage_output_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = MDSMixStage_output_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = MDSMixStage_output_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = MDSMixStage_output_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = MDSMixStage_output_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      AddRoundConstantStage_output_rValid <= 1'b0;
      AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      SBox5Stage_output_rValid <= 1'b0;
      SBox5Stage_output_m2sPipe_rValid <= 1'b0;
    end else begin
      if(AddRoundConstantStage_output_ready) begin
        AddRoundConstantStage_output_rValid <= AddRoundConstantStage_output_valid;
      end
      if(AddRoundConstantStage_output_m2sPipe_valid) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b1;
      end
      if(AddRoundConstantStage_output_m2sPipe_input_ready) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      end
      if(SBox5Stage_output_ready) begin
        SBox5Stage_output_rValid <= SBox5Stage_output_valid;
      end
      if(SBox5Stage_output_m2sPipe_valid) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b1;
      end
      if(SBox5Stage_output_m2sPipe_input_ready) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(AddRoundConstantStage_output_ready) begin
      AddRoundConstantStage_output_rData_round_index <= AddRoundConstantStage_output_payload_round_index;
      AddRoundConstantStage_output_rData_state_index <= AddRoundConstantStage_output_payload_state_index;
      AddRoundConstantStage_output_rData_state_size <= AddRoundConstantStage_output_payload_state_size;
      AddRoundConstantStage_output_rData_state_id <= AddRoundConstantStage_output_payload_state_id;
      AddRoundConstantStage_output_rData_state_element <= AddRoundConstantStage_output_payload_state_element;
    end
    if(AddRoundConstantStage_output_m2sPipe_ready) begin
      AddRoundConstantStage_output_m2sPipe_rData_round_index <= AddRoundConstantStage_output_m2sPipe_payload_round_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_index <= AddRoundConstantStage_output_m2sPipe_payload_state_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_size <= AddRoundConstantStage_output_m2sPipe_payload_state_size;
      AddRoundConstantStage_output_m2sPipe_rData_state_id <= AddRoundConstantStage_output_m2sPipe_payload_state_id;
      AddRoundConstantStage_output_m2sPipe_rData_state_element <= AddRoundConstantStage_output_m2sPipe_payload_state_element;
    end
    if(SBox5Stage_output_ready) begin
      SBox5Stage_output_rData_round_index <= SBox5Stage_output_payload_round_index;
      SBox5Stage_output_rData_state_index <= SBox5Stage_output_payload_state_index;
      SBox5Stage_output_rData_state_size <= SBox5Stage_output_payload_state_size;
      SBox5Stage_output_rData_state_id <= SBox5Stage_output_payload_state_id;
      SBox5Stage_output_rData_state_element <= SBox5Stage_output_payload_state_element;
    end
    if(SBox5Stage_output_m2sPipe_ready) begin
      SBox5Stage_output_m2sPipe_rData_round_index <= SBox5Stage_output_m2sPipe_payload_round_index;
      SBox5Stage_output_m2sPipe_rData_state_index <= SBox5Stage_output_m2sPipe_payload_state_index;
      SBox5Stage_output_m2sPipe_rData_state_size <= SBox5Stage_output_m2sPipe_payload_state_size;
      SBox5Stage_output_m2sPipe_rData_state_id <= SBox5Stage_output_m2sPipe_payload_state_id;
      SBox5Stage_output_m2sPipe_rData_state_element <= SBox5Stage_output_m2sPipe_payload_state_element;
    end
  end


endmodule

module PoseidonThread (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index;
  wire       [2:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index;
  wire       [5:0]    AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index;
  reg        [254:0]  AddRoundConstantStage_modAdder_op2_i;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
  wire       [254:0]  AddRoundConstantStage_modAdder_res_o;
  wire                SBox5Stage_SBox5Insts_0_io_input_ready;
  wire                SBox5Stage_SBox5Insts_0_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_0_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_0_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_1_io_input_ready;
  wire                SBox5Stage_SBox5Insts_1_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_1_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_1_io_output_payload_state_element;
  wire                SBox5Stage_SBox5Insts_2_io_input_ready;
  wire                SBox5Stage_SBox5Insts_2_io_output_valid;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_round_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_index;
  wire       [3:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_size;
  wire       [6:0]    SBox5Stage_SBox5Insts_2_io_output_payload_state_id;
  wire       [254:0]  SBox5Stage_SBox5Insts_2_io_output_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_0_payload_state_element;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_1_payload_state_element;
  wire                streamDemux_7_io_outputs_2_valid;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_7_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_7_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_7_io_outputs_2_payload_state_element;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [4:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_7_io_inputs_0_ready;
  wire                streamMux_7_io_inputs_1_ready;
  wire                streamMux_7_io_inputs_2_ready;
  wire                streamMux_7_io_output_valid;
  wire       [6:0]    streamMux_7_io_output_payload_round_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_index;
  wire       [3:0]    streamMux_7_io_output_payload_state_size;
  wire       [6:0]    streamMux_7_io_output_payload_state_id;
  wire       [254:0]  streamMux_7_io_output_payload_state_element;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_0_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_1_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_input_ready;
  wire                MDSMixStage_matrixMultiplierInsts_2_io_output_valid;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index;
  wire       [3:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size;
  wire       [6:0]    MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_input_ready;
  wire                streamDemux_8_io_outputs_0_valid;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_0_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_0_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_0_payload_state_element;
  wire                streamDemux_8_io_outputs_1_valid;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_1_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_1_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_1_payload_state_element;
  wire                streamDemux_8_io_outputs_2_valid;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_round_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_index;
  wire       [3:0]    streamDemux_8_io_outputs_2_payload_state_size;
  wire       [6:0]    streamDemux_8_io_outputs_2_payload_state_id;
  wire       [254:0]  streamDemux_8_io_outputs_2_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy;
  wire                streamMux_8_io_inputs_0_ready;
  wire                streamMux_8_io_inputs_1_ready;
  wire                streamMux_8_io_inputs_2_ready;
  wire                streamMux_8_io_output_valid;
  wire       [6:0]    streamMux_8_io_output_payload_round_index;
  wire       [3:0]    streamMux_8_io_output_payload_state_size;
  wire       [6:0]    streamMux_8_io_output_payload_state_id;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_0;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_1;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_2;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_3;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_4;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_5;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_6;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_7;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_8;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_9;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_10;
  wire       [254:0]  streamMux_8_io_output_payload_state_elements_11;
  wire       [2:0]    _zz__zz_SBox5Stage_DemuxSelect_1;
  wire       [2:0]    _zz__zz_MDSMixStage_DemuxSelect_1;
  wire                AddRoundConstantStage_output_valid;
  reg                 AddRoundConstantStage_output_ready;
  wire       [6:0]    AddRoundConstantStage_output_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_payload_state_id;
  reg        [254:0]  AddRoundConstantStage_output_payload_state_element;
  wire                when_PoseidonThread_l46;
  wire                AddRoundConstantStage_output_m2sPipe_valid;
  wire                AddRoundConstantStage_output_m2sPipe_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_payload_state_element;
  reg                 AddRoundConstantStage_output_rValid;
  reg        [6:0]    AddRoundConstantStage_output_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_rData_state_element;
  wire                when_Stream_l342;
  wire                AddRoundConstantStage_output_m2sPipe_input_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_ready;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    AddRoundConstantStage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  AddRoundConstantStage_output_m2sPipe_input_payload_state_element;
  reg                 AddRoundConstantStage_output_m2sPipe_rValid;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_round_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_index;
  reg        [3:0]    AddRoundConstantStage_output_m2sPipe_rData_state_size;
  reg        [6:0]    AddRoundConstantStage_output_m2sPipe_rData_state_id;
  reg        [254:0]  AddRoundConstantStage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect;
  wire       [2:0]    _zz_SBox5Stage_DemuxSelect_1;
  wire                _zz_SBox5Stage_DemuxSelect_2;
  wire                _zz_SBox5Stage_DemuxSelect_3;
  wire       [1:0]    SBox5Stage_DemuxSelect;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_SBox5Stage_output_valid;
  wire                _zz_io_pop_ready;
  wire                SBox5Stage_output_valid;
  reg                 SBox5Stage_output_ready;
  wire       [6:0]    SBox5Stage_output_payload_round_index;
  wire       [3:0]    SBox5Stage_output_payload_state_index;
  wire       [3:0]    SBox5Stage_output_payload_state_size;
  wire       [6:0]    SBox5Stage_output_payload_state_id;
  wire       [254:0]  SBox5Stage_output_payload_state_element;
  wire                SBox5Stage_output_m2sPipe_valid;
  wire                SBox5Stage_output_m2sPipe_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_payload_state_element;
  reg                 SBox5Stage_output_rValid;
  reg        [6:0]    SBox5Stage_output_rData_round_index;
  reg        [3:0]    SBox5Stage_output_rData_state_index;
  reg        [3:0]    SBox5Stage_output_rData_state_size;
  reg        [6:0]    SBox5Stage_output_rData_state_id;
  reg        [254:0]  SBox5Stage_output_rData_state_element;
  wire                when_Stream_l342_1;
  wire                SBox5Stage_output_m2sPipe_input_valid;
  wire                SBox5Stage_output_m2sPipe_input_ready;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_round_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_index;
  wire       [3:0]    SBox5Stage_output_m2sPipe_input_payload_state_size;
  wire       [6:0]    SBox5Stage_output_m2sPipe_input_payload_state_id;
  wire       [254:0]  SBox5Stage_output_m2sPipe_input_payload_state_element;
  reg                 SBox5Stage_output_m2sPipe_rValid;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_round_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_index;
  reg        [3:0]    SBox5Stage_output_m2sPipe_rData_state_size;
  reg        [6:0]    SBox5Stage_output_m2sPipe_rData_state_id;
  reg        [254:0]  SBox5Stage_output_m2sPipe_rData_state_element;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect;
  wire       [2:0]    _zz_MDSMixStage_DemuxSelect_1;
  wire                _zz_MDSMixStage_DemuxSelect_2;
  wire                _zz_MDSMixStage_DemuxSelect_3;
  wire       [1:0]    MDSMixStage_DemuxSelect;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid;
  wire                SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready;
  wire       [1:0]    SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload;
  wire                _zz_MDSMixStage_output_valid;
  wire                _zz_io_pop_ready_1;
  wire                MDSMixStage_output_valid;
  wire                MDSMixStage_output_ready;
  wire       [6:0]    MDSMixStage_output_payload_round_index;
  wire       [3:0]    MDSMixStage_output_payload_state_size;
  wire       [6:0]    MDSMixStage_output_payload_state_id;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_0;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_1;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_2;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_3;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_4;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_5;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_6;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_7;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_8;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_9;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_10;
  wire       [254:0]  MDSMixStage_output_payload_state_elements_11;

  assign _zz__zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect - 3'b001);
  assign _zz__zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect - 3'b001);
  RoundConstants AddRoundConstantStage_roundConstants_t3 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_1 AddRoundConstantStage_roundConstants_t5 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data         ), //o
    .io_read_ports_0_t_index        (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index      ), //i
    .io_read_ports_0_round_index    (AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index  )  //i
  );
  RoundConstants_2 AddRoundConstantStage_roundConstants_t9 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                  ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                  )  //i
  );
  RoundConstants_3 AddRoundConstantStage_roundConstants_t12 (
    .io_read_ports_0_data           (AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data  ), //o
    .io_read_ports_0_t_index        (io_input_payload_state_index                                   ), //i
    .io_read_ports_0_round_index    (io_input_payload_round_index                                   )  //i
  );
  ModAdder AddRoundConstantStage_modAdder (
    .op1_i    (io_input_payload_state_element        ), //i
    .op2_i    (AddRoundConstantStage_modAdder_op2_i  ), //i
    .res_o    (AddRoundConstantStage_modAdder_res_o  )  //o
  );
  SBox5 SBox5Stage_SBox5Insts_0 (
    .io_input_valid                     (streamDemux_7_io_outputs_0_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_0_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_0_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_0_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_0_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_0_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_0_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_0_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_1 (
    .io_input_valid                     (streamDemux_7_io_outputs_1_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_1_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_1_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_1_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_1_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_1_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_1_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_1_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  SBox5 SBox5Stage_SBox5Insts_2 (
    .io_input_valid                     (streamDemux_7_io_outputs_2_valid                         ), //i
    .io_input_ready                     (SBox5Stage_SBox5Insts_2_io_input_ready                   ), //o
    .io_input_payload_round_index       (streamDemux_7_io_outputs_2_payload_round_index           ), //i
    .io_input_payload_state_index       (streamDemux_7_io_outputs_2_payload_state_index           ), //i
    .io_input_payload_state_size        (streamDemux_7_io_outputs_2_payload_state_size            ), //i
    .io_input_payload_state_id          (streamDemux_7_io_outputs_2_payload_state_id              ), //i
    .io_input_payload_state_element     (streamDemux_7_io_outputs_2_payload_state_element         ), //i
    .io_output_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                  ), //o
    .io_output_ready                    (streamMux_7_io_inputs_2_ready                            ), //i
    .io_output_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index    ), //o
    .io_output_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index    ), //o
    .io_output_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size     ), //o
    .io_output_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id       ), //o
    .io_output_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element  ), //o
    .reset                              (reset                                                    ), //i
    .clk                                (clk                                                      )  //i
  );
  StreamFork_10 AddRoundConstantStage_output_m2sPipe_input_fork (
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_7_io_input_ready                                                        ), //i
    .io_outputs_0_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_7 (
    .io_select                             (SBox5Stage_DemuxSelect                                                              ), //i
    .io_input_valid                        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_7_io_input_ready                                                        ), //o
    .io_input_payload_round_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_7_io_outputs_0_valid                                                    ), //o
    .io_outputs_0_ready                    (SBox5Stage_SBox5Insts_0_io_input_ready                                              ), //i
    .io_outputs_0_payload_round_index      (streamDemux_7_io_outputs_0_payload_round_index                                      ), //o
    .io_outputs_0_payload_state_index      (streamDemux_7_io_outputs_0_payload_state_index                                      ), //o
    .io_outputs_0_payload_state_size       (streamDemux_7_io_outputs_0_payload_state_size                                       ), //o
    .io_outputs_0_payload_state_id         (streamDemux_7_io_outputs_0_payload_state_id                                         ), //o
    .io_outputs_0_payload_state_element    (streamDemux_7_io_outputs_0_payload_state_element                                    ), //o
    .io_outputs_1_valid                    (streamDemux_7_io_outputs_1_valid                                                    ), //o
    .io_outputs_1_ready                    (SBox5Stage_SBox5Insts_1_io_input_ready                                              ), //i
    .io_outputs_1_payload_round_index      (streamDemux_7_io_outputs_1_payload_round_index                                      ), //o
    .io_outputs_1_payload_state_index      (streamDemux_7_io_outputs_1_payload_state_index                                      ), //o
    .io_outputs_1_payload_state_size       (streamDemux_7_io_outputs_1_payload_state_size                                       ), //o
    .io_outputs_1_payload_state_id         (streamDemux_7_io_outputs_1_payload_state_id                                         ), //o
    .io_outputs_1_payload_state_element    (streamDemux_7_io_outputs_1_payload_state_element                                    ), //o
    .io_outputs_2_valid                    (streamDemux_7_io_outputs_2_valid                                                    ), //o
    .io_outputs_2_ready                    (SBox5Stage_SBox5Insts_2_io_input_ready                                              ), //i
    .io_outputs_2_payload_round_index      (streamDemux_7_io_outputs_2_payload_round_index                                      ), //o
    .io_outputs_2_payload_state_index      (streamDemux_7_io_outputs_2_payload_state_index                                      ), //o
    .io_outputs_2_payload_state_size       (streamDemux_7_io_outputs_2_payload_state_size                                       ), //o
    .io_outputs_2_payload_state_id         (streamDemux_7_io_outputs_2_payload_state_id                                         ), //o
    .io_outputs_2_payload_state_element    (streamDemux_7_io_outputs_2_payload_state_element                                    )  //o
  );
  StreamFifoLowLatency AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready                                                                             ), //i
    .io_pop_payload     (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                                         ), //i
    .io_occupancy       (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                                          ), //i
    .reset              (reset                                                                                        )  //i
  );
  StreamMux streamMux_7 (
    .io_select                            (AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                    (SBox5Stage_SBox5Insts_0_io_output_valid                                                      ), //i
    .io_inputs_0_ready                    (streamMux_7_io_inputs_0_ready                                                                ), //o
    .io_inputs_0_payload_round_index      (SBox5Stage_SBox5Insts_0_io_output_payload_round_index                                        ), //i
    .io_inputs_0_payload_state_index      (SBox5Stage_SBox5Insts_0_io_output_payload_state_index                                        ), //i
    .io_inputs_0_payload_state_size       (SBox5Stage_SBox5Insts_0_io_output_payload_state_size                                         ), //i
    .io_inputs_0_payload_state_id         (SBox5Stage_SBox5Insts_0_io_output_payload_state_id                                           ), //i
    .io_inputs_0_payload_state_element    (SBox5Stage_SBox5Insts_0_io_output_payload_state_element                                      ), //i
    .io_inputs_1_valid                    (SBox5Stage_SBox5Insts_1_io_output_valid                                                      ), //i
    .io_inputs_1_ready                    (streamMux_7_io_inputs_1_ready                                                                ), //o
    .io_inputs_1_payload_round_index      (SBox5Stage_SBox5Insts_1_io_output_payload_round_index                                        ), //i
    .io_inputs_1_payload_state_index      (SBox5Stage_SBox5Insts_1_io_output_payload_state_index                                        ), //i
    .io_inputs_1_payload_state_size       (SBox5Stage_SBox5Insts_1_io_output_payload_state_size                                         ), //i
    .io_inputs_1_payload_state_id         (SBox5Stage_SBox5Insts_1_io_output_payload_state_id                                           ), //i
    .io_inputs_1_payload_state_element    (SBox5Stage_SBox5Insts_1_io_output_payload_state_element                                      ), //i
    .io_inputs_2_valid                    (SBox5Stage_SBox5Insts_2_io_output_valid                                                      ), //i
    .io_inputs_2_ready                    (streamMux_7_io_inputs_2_ready                                                                ), //o
    .io_inputs_2_payload_round_index      (SBox5Stage_SBox5Insts_2_io_output_payload_round_index                                        ), //i
    .io_inputs_2_payload_state_index      (SBox5Stage_SBox5Insts_2_io_output_payload_state_index                                        ), //i
    .io_inputs_2_payload_state_size       (SBox5Stage_SBox5Insts_2_io_output_payload_state_size                                         ), //i
    .io_inputs_2_payload_state_id         (SBox5Stage_SBox5Insts_2_io_output_payload_state_id                                           ), //i
    .io_inputs_2_payload_state_element    (SBox5Stage_SBox5Insts_2_io_output_payload_state_element                                      ), //i
    .io_output_valid                      (streamMux_7_io_output_valid                                                                  ), //o
    .io_output_ready                      (_zz_io_pop_ready                                                                             ), //i
    .io_output_payload_round_index        (streamMux_7_io_output_payload_round_index                                                    ), //o
    .io_output_payload_state_index        (streamMux_7_io_output_payload_state_index                                                    ), //o
    .io_output_payload_state_size         (streamMux_7_io_output_payload_state_size                                                     ), //o
    .io_output_payload_state_id           (streamMux_7_io_output_payload_state_id                                                       ), //o
    .io_output_payload_state_element      (streamMux_7_io_output_payload_state_element                                                  )  //o
  );
  MDSMatrixMultiplier MDSMixStage_matrixMultiplierInsts_0 (
    .io_input_valid                         (streamDemux_8_io_outputs_0_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_0_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_0_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_0_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_0_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_0_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_0_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_1 MDSMixStage_matrixMultiplierInsts_1 (
    .io_input_valid                         (streamDemux_8_io_outputs_1_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_1_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_1_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_1_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_1_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_1_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_1_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  MDSMatrixMultiplier_2 MDSMixStage_matrixMultiplierInsts_2 (
    .io_input_valid                         (streamDemux_8_io_outputs_2_valid                                         ), //i
    .io_input_ready                         (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //o
    .io_input_payload_round_index           (streamDemux_8_io_outputs_2_payload_round_index                           ), //i
    .io_input_payload_state_index           (streamDemux_8_io_outputs_2_payload_state_index                           ), //i
    .io_input_payload_state_size            (streamDemux_8_io_outputs_2_payload_state_size                            ), //i
    .io_input_payload_state_id              (streamDemux_8_io_outputs_2_payload_state_id                              ), //i
    .io_input_payload_state_element         (streamDemux_8_io_outputs_2_payload_state_element                         ), //i
    .io_output_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                      ), //o
    .io_output_ready                        (streamMux_8_io_inputs_2_ready                                            ), //i
    .io_output_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index        ), //o
    .io_output_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size         ), //o
    .io_output_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id           ), //o
    .io_output_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0   ), //o
    .io_output_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1   ), //o
    .io_output_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2   ), //o
    .io_output_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3   ), //o
    .io_output_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4   ), //o
    .io_output_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5   ), //o
    .io_output_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6   ), //o
    .io_output_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7   ), //o
    .io_output_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8   ), //o
    .io_output_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9   ), //o
    .io_output_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10  ), //o
    .io_output_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11  ), //o
    .reset                                  (reset                                                                    ), //i
    .clk                                    (clk                                                                      )  //i
  );
  StreamFork_10 SBox5Stage_output_m2sPipe_input_fork (
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_valid                                    ), //i
    .io_input_ready                        (SBox5Stage_output_m2sPipe_input_fork_io_input_ready                      ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_payload_round_index                      ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_payload_state_index                      ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_payload_state_size                       ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_payload_state_id                         ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_payload_state_element                    ), //i
    .io_outputs_0_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //o
    .io_outputs_0_ready                    (streamDemux_8_io_input_ready                                             ), //i
    .io_outputs_0_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //o
    .io_outputs_0_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //o
    .io_outputs_0_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //o
    .io_outputs_0_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //o
    .io_outputs_0_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //o
    .io_outputs_1_valid                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid                  ), //o
    .io_outputs_1_ready                    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready       ), //i
    .io_outputs_1_payload_round_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_round_index    ), //o
    .io_outputs_1_payload_state_index      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_index    ), //o
    .io_outputs_1_payload_state_size       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_size     ), //o
    .io_outputs_1_payload_state_id         (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_id       ), //o
    .io_outputs_1_payload_state_element    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_payload_state_element  )  //o
  );
  StreamDemux streamDemux_8 (
    .io_select                             (MDSMixStage_DemuxSelect                                                  ), //i
    .io_input_valid                        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_valid                  ), //i
    .io_input_ready                        (streamDemux_8_io_input_ready                                             ), //o
    .io_input_payload_round_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_round_index    ), //i
    .io_input_payload_state_index          (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_index    ), //i
    .io_input_payload_state_size           (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_size     ), //i
    .io_input_payload_state_id             (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_id       ), //i
    .io_input_payload_state_element        (SBox5Stage_output_m2sPipe_input_fork_io_outputs_0_payload_state_element  ), //i
    .io_outputs_0_valid                    (streamDemux_8_io_outputs_0_valid                                         ), //o
    .io_outputs_0_ready                    (MDSMixStage_matrixMultiplierInsts_0_io_input_ready                       ), //i
    .io_outputs_0_payload_round_index      (streamDemux_8_io_outputs_0_payload_round_index                           ), //o
    .io_outputs_0_payload_state_index      (streamDemux_8_io_outputs_0_payload_state_index                           ), //o
    .io_outputs_0_payload_state_size       (streamDemux_8_io_outputs_0_payload_state_size                            ), //o
    .io_outputs_0_payload_state_id         (streamDemux_8_io_outputs_0_payload_state_id                              ), //o
    .io_outputs_0_payload_state_element    (streamDemux_8_io_outputs_0_payload_state_element                         ), //o
    .io_outputs_1_valid                    (streamDemux_8_io_outputs_1_valid                                         ), //o
    .io_outputs_1_ready                    (MDSMixStage_matrixMultiplierInsts_1_io_input_ready                       ), //i
    .io_outputs_1_payload_round_index      (streamDemux_8_io_outputs_1_payload_round_index                           ), //o
    .io_outputs_1_payload_state_index      (streamDemux_8_io_outputs_1_payload_state_index                           ), //o
    .io_outputs_1_payload_state_size       (streamDemux_8_io_outputs_1_payload_state_size                            ), //o
    .io_outputs_1_payload_state_id         (streamDemux_8_io_outputs_1_payload_state_id                              ), //o
    .io_outputs_1_payload_state_element    (streamDemux_8_io_outputs_1_payload_state_element                         ), //o
    .io_outputs_2_valid                    (streamDemux_8_io_outputs_2_valid                                         ), //o
    .io_outputs_2_ready                    (MDSMixStage_matrixMultiplierInsts_2_io_input_ready                       ), //i
    .io_outputs_2_payload_round_index      (streamDemux_8_io_outputs_2_payload_round_index                           ), //o
    .io_outputs_2_payload_state_index      (streamDemux_8_io_outputs_2_payload_state_index                           ), //o
    .io_outputs_2_payload_state_size       (streamDemux_8_io_outputs_2_payload_state_size                            ), //o
    .io_outputs_2_payload_state_id         (streamDemux_8_io_outputs_2_payload_state_id                              ), //o
    .io_outputs_2_payload_state_element    (streamDemux_8_io_outputs_2_payload_state_element                         )  //o
  );
  StreamFifoLowLatency_1 SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo (
    .io_push_valid      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid                ), //i
    .io_push_ready      (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready   ), //o
    .io_push_payload    (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload              ), //i
    .io_pop_valid       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid    ), //o
    .io_pop_ready       (_zz_io_pop_ready_1                                                                ), //i
    .io_pop_payload     (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //o
    .io_flush           (1'b0                                                                              ), //i
    .io_occupancy       (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_occupancy    ), //o
    .clk                (clk                                                                               ), //i
    .reset              (reset                                                                             )  //i
  );
  StreamMux_1 streamMux_8 (
    .io_select                                (SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_payload  ), //i
    .io_inputs_0_valid                        (MDSMixStage_matrixMultiplierInsts_0_io_output_valid                               ), //i
    .io_inputs_0_ready                        (streamMux_8_io_inputs_0_ready                                                     ), //o
    .io_inputs_0_payload_round_index          (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_round_index                 ), //i
    .io_inputs_0_payload_state_size           (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_size                  ), //i
    .io_inputs_0_payload_state_id             (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_id                    ), //i
    .io_inputs_0_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_0            ), //i
    .io_inputs_0_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_1            ), //i
    .io_inputs_0_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_2            ), //i
    .io_inputs_0_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_3            ), //i
    .io_inputs_0_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_4            ), //i
    .io_inputs_0_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_5            ), //i
    .io_inputs_0_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_6            ), //i
    .io_inputs_0_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_7            ), //i
    .io_inputs_0_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_8            ), //i
    .io_inputs_0_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_9            ), //i
    .io_inputs_0_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_10           ), //i
    .io_inputs_0_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_0_io_output_payload_state_elements_11           ), //i
    .io_inputs_1_valid                        (MDSMixStage_matrixMultiplierInsts_1_io_output_valid                               ), //i
    .io_inputs_1_ready                        (streamMux_8_io_inputs_1_ready                                                     ), //o
    .io_inputs_1_payload_round_index          (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_round_index                 ), //i
    .io_inputs_1_payload_state_size           (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_size                  ), //i
    .io_inputs_1_payload_state_id             (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_id                    ), //i
    .io_inputs_1_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_0            ), //i
    .io_inputs_1_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_1            ), //i
    .io_inputs_1_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_2            ), //i
    .io_inputs_1_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_3            ), //i
    .io_inputs_1_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_4            ), //i
    .io_inputs_1_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_5            ), //i
    .io_inputs_1_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_6            ), //i
    .io_inputs_1_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_7            ), //i
    .io_inputs_1_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_8            ), //i
    .io_inputs_1_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_9            ), //i
    .io_inputs_1_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_10           ), //i
    .io_inputs_1_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_1_io_output_payload_state_elements_11           ), //i
    .io_inputs_2_valid                        (MDSMixStage_matrixMultiplierInsts_2_io_output_valid                               ), //i
    .io_inputs_2_ready                        (streamMux_8_io_inputs_2_ready                                                     ), //o
    .io_inputs_2_payload_round_index          (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_round_index                 ), //i
    .io_inputs_2_payload_state_size           (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_size                  ), //i
    .io_inputs_2_payload_state_id             (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_id                    ), //i
    .io_inputs_2_payload_state_elements_0     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_0            ), //i
    .io_inputs_2_payload_state_elements_1     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_1            ), //i
    .io_inputs_2_payload_state_elements_2     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_2            ), //i
    .io_inputs_2_payload_state_elements_3     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_3            ), //i
    .io_inputs_2_payload_state_elements_4     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_4            ), //i
    .io_inputs_2_payload_state_elements_5     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_5            ), //i
    .io_inputs_2_payload_state_elements_6     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_6            ), //i
    .io_inputs_2_payload_state_elements_7     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_7            ), //i
    .io_inputs_2_payload_state_elements_8     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_8            ), //i
    .io_inputs_2_payload_state_elements_9     (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_9            ), //i
    .io_inputs_2_payload_state_elements_10    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_10           ), //i
    .io_inputs_2_payload_state_elements_11    (MDSMixStage_matrixMultiplierInsts_2_io_output_payload_state_elements_11           ), //i
    .io_output_valid                          (streamMux_8_io_output_valid                                                       ), //o
    .io_output_ready                          (_zz_io_pop_ready_1                                                                ), //i
    .io_output_payload_round_index            (streamMux_8_io_output_payload_round_index                                         ), //o
    .io_output_payload_state_size             (streamMux_8_io_output_payload_state_size                                          ), //o
    .io_output_payload_state_id               (streamMux_8_io_output_payload_state_id                                            ), //o
    .io_output_payload_state_elements_0       (streamMux_8_io_output_payload_state_elements_0                                    ), //o
    .io_output_payload_state_elements_1       (streamMux_8_io_output_payload_state_elements_1                                    ), //o
    .io_output_payload_state_elements_2       (streamMux_8_io_output_payload_state_elements_2                                    ), //o
    .io_output_payload_state_elements_3       (streamMux_8_io_output_payload_state_elements_3                                    ), //o
    .io_output_payload_state_elements_4       (streamMux_8_io_output_payload_state_elements_4                                    ), //o
    .io_output_payload_state_elements_5       (streamMux_8_io_output_payload_state_elements_5                                    ), //o
    .io_output_payload_state_elements_6       (streamMux_8_io_output_payload_state_elements_6                                    ), //o
    .io_output_payload_state_elements_7       (streamMux_8_io_output_payload_state_elements_7                                    ), //o
    .io_output_payload_state_elements_8       (streamMux_8_io_output_payload_state_elements_8                                    ), //o
    .io_output_payload_state_elements_9       (streamMux_8_io_output_payload_state_elements_9                                    ), //o
    .io_output_payload_state_elements_10      (streamMux_8_io_output_payload_state_elements_10                                   ), //o
    .io_output_payload_state_elements_11      (streamMux_8_io_output_payload_state_elements_11                                   )  //o
  );
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_t_index = io_input_payload_state_index[1:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_t_index = io_input_payload_state_index[2:0];
  assign AddRoundConstantStage_roundConstants_t3_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  assign AddRoundConstantStage_roundConstants_t5_io_read_ports_0_round_index = io_input_payload_round_index[5:0];
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t3_io_read_ports_0_data;
      end
      4'b0101 : begin
        if(when_PoseidonThread_l46) begin
          AddRoundConstantStage_modAdder_op2_i = 255'h0;
        end else begin
          AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t5_io_read_ports_0_data;
        end
      end
      4'b1001 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t9_io_read_ports_0_data;
      end
      4'b1100 : begin
        AddRoundConstantStage_modAdder_op2_i = AddRoundConstantStage_roundConstants_t12_io_read_ports_0_data;
      end
      default : begin
        AddRoundConstantStage_modAdder_op2_i = 255'h0;
      end
    endcase
  end

  assign when_PoseidonThread_l46 = (io_input_payload_state_index == 4'b0101);
  assign AddRoundConstantStage_output_valid = io_input_valid;
  assign io_input_ready = AddRoundConstantStage_output_ready;
  assign AddRoundConstantStage_output_payload_round_index = io_input_payload_round_index;
  assign AddRoundConstantStage_output_payload_state_index = io_input_payload_state_index;
  assign AddRoundConstantStage_output_payload_state_size = io_input_payload_state_size;
  assign AddRoundConstantStage_output_payload_state_id = io_input_payload_state_id;
  always @(*) begin
    AddRoundConstantStage_output_payload_state_element = io_input_payload_state_element;
    AddRoundConstantStage_output_payload_state_element = AddRoundConstantStage_modAdder_res_o;
  end

  always @(*) begin
    AddRoundConstantStage_output_ready = AddRoundConstantStage_output_m2sPipe_ready;
    if(when_Stream_l342) begin
      AddRoundConstantStage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! AddRoundConstantStage_output_m2sPipe_valid);
  assign AddRoundConstantStage_output_m2sPipe_valid = AddRoundConstantStage_output_rValid;
  assign AddRoundConstantStage_output_m2sPipe_payload_round_index = AddRoundConstantStage_output_rData_round_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_index = AddRoundConstantStage_output_rData_state_index;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_size = AddRoundConstantStage_output_rData_state_size;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_id = AddRoundConstantStage_output_rData_state_id;
  assign AddRoundConstantStage_output_m2sPipe_payload_state_element = AddRoundConstantStage_output_rData_state_element;
  assign AddRoundConstantStage_output_m2sPipe_ready = (! AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_valid = (AddRoundConstantStage_output_m2sPipe_valid || AddRoundConstantStage_output_m2sPipe_rValid);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_round_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_round_index : AddRoundConstantStage_output_m2sPipe_payload_round_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_index = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_index : AddRoundConstantStage_output_m2sPipe_payload_state_index);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_size = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_size : AddRoundConstantStage_output_m2sPipe_payload_state_size);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_id = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_id : AddRoundConstantStage_output_m2sPipe_payload_state_id);
  assign AddRoundConstantStage_output_m2sPipe_input_payload_state_element = (AddRoundConstantStage_output_m2sPipe_rValid ? AddRoundConstantStage_output_m2sPipe_rData_state_element : AddRoundConstantStage_output_m2sPipe_payload_state_element);
  assign AddRoundConstantStage_output_m2sPipe_input_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_SBox5Stage_DemuxSelect = {SBox5Stage_SBox5Insts_2_io_input_ready,{SBox5Stage_SBox5Insts_1_io_input_ready,SBox5Stage_SBox5Insts_0_io_input_ready}};
  assign _zz_SBox5Stage_DemuxSelect_1 = (_zz_SBox5Stage_DemuxSelect & (~ _zz__zz_SBox5Stage_DemuxSelect_1));
  assign _zz_SBox5Stage_DemuxSelect_2 = _zz_SBox5Stage_DemuxSelect_1[1];
  assign _zz_SBox5Stage_DemuxSelect_3 = _zz_SBox5Stage_DemuxSelect_1[2];
  assign SBox5Stage_DemuxSelect = {_zz_SBox5Stage_DemuxSelect_3,_zz_SBox5Stage_DemuxSelect_2};
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = SBox5Stage_DemuxSelect;
  assign AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready = (_zz_SBox5Stage_output_valid && SBox5Stage_output_ready);
  assign _zz_SBox5Stage_output_valid = (streamMux_7_io_output_valid && AddRoundConstantStage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign SBox5Stage_output_valid = _zz_SBox5Stage_output_valid;
  assign SBox5Stage_output_payload_round_index = streamMux_7_io_output_payload_round_index;
  assign SBox5Stage_output_payload_state_index = streamMux_7_io_output_payload_state_index;
  assign SBox5Stage_output_payload_state_size = streamMux_7_io_output_payload_state_size;
  assign SBox5Stage_output_payload_state_id = streamMux_7_io_output_payload_state_id;
  assign SBox5Stage_output_payload_state_element = streamMux_7_io_output_payload_state_element;
  always @(*) begin
    SBox5Stage_output_ready = SBox5Stage_output_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      SBox5Stage_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! SBox5Stage_output_m2sPipe_valid);
  assign SBox5Stage_output_m2sPipe_valid = SBox5Stage_output_rValid;
  assign SBox5Stage_output_m2sPipe_payload_round_index = SBox5Stage_output_rData_round_index;
  assign SBox5Stage_output_m2sPipe_payload_state_index = SBox5Stage_output_rData_state_index;
  assign SBox5Stage_output_m2sPipe_payload_state_size = SBox5Stage_output_rData_state_size;
  assign SBox5Stage_output_m2sPipe_payload_state_id = SBox5Stage_output_rData_state_id;
  assign SBox5Stage_output_m2sPipe_payload_state_element = SBox5Stage_output_rData_state_element;
  assign SBox5Stage_output_m2sPipe_ready = (! SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_valid = (SBox5Stage_output_m2sPipe_valid || SBox5Stage_output_m2sPipe_rValid);
  assign SBox5Stage_output_m2sPipe_input_payload_round_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_round_index : SBox5Stage_output_m2sPipe_payload_round_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_index = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_index : SBox5Stage_output_m2sPipe_payload_state_index);
  assign SBox5Stage_output_m2sPipe_input_payload_state_size = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_size : SBox5Stage_output_m2sPipe_payload_state_size);
  assign SBox5Stage_output_m2sPipe_input_payload_state_id = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_id : SBox5Stage_output_m2sPipe_payload_state_id);
  assign SBox5Stage_output_m2sPipe_input_payload_state_element = (SBox5Stage_output_m2sPipe_rValid ? SBox5Stage_output_m2sPipe_rData_state_element : SBox5Stage_output_m2sPipe_payload_state_element);
  assign SBox5Stage_output_m2sPipe_input_ready = SBox5Stage_output_m2sPipe_input_fork_io_input_ready;
  assign _zz_MDSMixStage_DemuxSelect = {MDSMixStage_matrixMultiplierInsts_2_io_input_ready,{MDSMixStage_matrixMultiplierInsts_1_io_input_ready,MDSMixStage_matrixMultiplierInsts_0_io_input_ready}};
  assign _zz_MDSMixStage_DemuxSelect_1 = (_zz_MDSMixStage_DemuxSelect & (~ _zz__zz_MDSMixStage_DemuxSelect_1));
  assign _zz_MDSMixStage_DemuxSelect_2 = _zz_MDSMixStage_DemuxSelect_1[1];
  assign _zz_MDSMixStage_DemuxSelect_3 = _zz_MDSMixStage_DemuxSelect_1[2];
  assign MDSMixStage_DemuxSelect = {_zz_MDSMixStage_DemuxSelect_3,_zz_MDSMixStage_DemuxSelect_2};
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_valid = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_valid;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_payload = MDSMixStage_DemuxSelect;
  assign SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_ready = SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_push_ready;
  assign _zz_io_pop_ready_1 = (_zz_MDSMixStage_output_valid && MDSMixStage_output_ready);
  assign _zz_MDSMixStage_output_valid = (streamMux_8_io_output_valid && SBox5Stage_output_m2sPipe_input_fork_io_outputs_1_translated_fifo_io_pop_valid);
  assign MDSMixStage_output_valid = _zz_MDSMixStage_output_valid;
  assign MDSMixStage_output_payload_round_index = streamMux_8_io_output_payload_round_index;
  assign MDSMixStage_output_payload_state_size = streamMux_8_io_output_payload_state_size;
  assign MDSMixStage_output_payload_state_id = streamMux_8_io_output_payload_state_id;
  assign MDSMixStage_output_payload_state_elements_0 = streamMux_8_io_output_payload_state_elements_0;
  assign MDSMixStage_output_payload_state_elements_1 = streamMux_8_io_output_payload_state_elements_1;
  assign MDSMixStage_output_payload_state_elements_2 = streamMux_8_io_output_payload_state_elements_2;
  assign MDSMixStage_output_payload_state_elements_3 = streamMux_8_io_output_payload_state_elements_3;
  assign MDSMixStage_output_payload_state_elements_4 = streamMux_8_io_output_payload_state_elements_4;
  assign MDSMixStage_output_payload_state_elements_5 = streamMux_8_io_output_payload_state_elements_5;
  assign MDSMixStage_output_payload_state_elements_6 = streamMux_8_io_output_payload_state_elements_6;
  assign MDSMixStage_output_payload_state_elements_7 = streamMux_8_io_output_payload_state_elements_7;
  assign MDSMixStage_output_payload_state_elements_8 = streamMux_8_io_output_payload_state_elements_8;
  assign MDSMixStage_output_payload_state_elements_9 = streamMux_8_io_output_payload_state_elements_9;
  assign MDSMixStage_output_payload_state_elements_10 = streamMux_8_io_output_payload_state_elements_10;
  assign MDSMixStage_output_payload_state_elements_11 = streamMux_8_io_output_payload_state_elements_11;
  assign io_output_valid = MDSMixStage_output_valid;
  assign MDSMixStage_output_ready = io_output_ready;
  assign io_output_payload_round_index = MDSMixStage_output_payload_round_index;
  assign io_output_payload_state_size = MDSMixStage_output_payload_state_size;
  assign io_output_payload_state_id = MDSMixStage_output_payload_state_id;
  assign io_output_payload_state_elements_0 = MDSMixStage_output_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = MDSMixStage_output_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = MDSMixStage_output_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = MDSMixStage_output_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = MDSMixStage_output_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = MDSMixStage_output_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = MDSMixStage_output_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = MDSMixStage_output_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = MDSMixStage_output_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = MDSMixStage_output_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = MDSMixStage_output_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = MDSMixStage_output_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      AddRoundConstantStage_output_rValid <= 1'b0;
      AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      SBox5Stage_output_rValid <= 1'b0;
      SBox5Stage_output_m2sPipe_rValid <= 1'b0;
    end else begin
      if(AddRoundConstantStage_output_ready) begin
        AddRoundConstantStage_output_rValid <= AddRoundConstantStage_output_valid;
      end
      if(AddRoundConstantStage_output_m2sPipe_valid) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b1;
      end
      if(AddRoundConstantStage_output_m2sPipe_input_ready) begin
        AddRoundConstantStage_output_m2sPipe_rValid <= 1'b0;
      end
      if(SBox5Stage_output_ready) begin
        SBox5Stage_output_rValid <= SBox5Stage_output_valid;
      end
      if(SBox5Stage_output_m2sPipe_valid) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b1;
      end
      if(SBox5Stage_output_m2sPipe_input_ready) begin
        SBox5Stage_output_m2sPipe_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(AddRoundConstantStage_output_ready) begin
      AddRoundConstantStage_output_rData_round_index <= AddRoundConstantStage_output_payload_round_index;
      AddRoundConstantStage_output_rData_state_index <= AddRoundConstantStage_output_payload_state_index;
      AddRoundConstantStage_output_rData_state_size <= AddRoundConstantStage_output_payload_state_size;
      AddRoundConstantStage_output_rData_state_id <= AddRoundConstantStage_output_payload_state_id;
      AddRoundConstantStage_output_rData_state_element <= AddRoundConstantStage_output_payload_state_element;
    end
    if(AddRoundConstantStage_output_m2sPipe_ready) begin
      AddRoundConstantStage_output_m2sPipe_rData_round_index <= AddRoundConstantStage_output_m2sPipe_payload_round_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_index <= AddRoundConstantStage_output_m2sPipe_payload_state_index;
      AddRoundConstantStage_output_m2sPipe_rData_state_size <= AddRoundConstantStage_output_m2sPipe_payload_state_size;
      AddRoundConstantStage_output_m2sPipe_rData_state_id <= AddRoundConstantStage_output_m2sPipe_payload_state_id;
      AddRoundConstantStage_output_m2sPipe_rData_state_element <= AddRoundConstantStage_output_m2sPipe_payload_state_element;
    end
    if(SBox5Stage_output_ready) begin
      SBox5Stage_output_rData_round_index <= SBox5Stage_output_payload_round_index;
      SBox5Stage_output_rData_state_index <= SBox5Stage_output_payload_state_index;
      SBox5Stage_output_rData_state_size <= SBox5Stage_output_payload_state_size;
      SBox5Stage_output_rData_state_id <= SBox5Stage_output_payload_state_id;
      SBox5Stage_output_rData_state_element <= SBox5Stage_output_payload_state_element;
    end
    if(SBox5Stage_output_m2sPipe_ready) begin
      SBox5Stage_output_m2sPipe_rData_round_index <= SBox5Stage_output_m2sPipe_payload_round_index;
      SBox5Stage_output_m2sPipe_rData_state_index <= SBox5Stage_output_m2sPipe_payload_state_index;
      SBox5Stage_output_m2sPipe_rData_state_size <= SBox5Stage_output_m2sPipe_payload_state_size;
      SBox5Stage_output_m2sPipe_rData_state_id <= SBox5Stage_output_m2sPipe_payload_state_id;
      SBox5Stage_output_m2sPipe_rData_state_element <= SBox5Stage_output_m2sPipe_payload_state_element;
    end
  end


endmodule

module MDSMatrixAdders (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [6:0]    io_inputs_0_payload_round_index,
  input      [3:0]    io_inputs_0_payload_state_size,
  input      [6:0]    io_inputs_0_payload_state_id,
  input      [254:0]  io_inputs_0_payload_state_elements_0,
  input      [254:0]  io_inputs_0_payload_state_elements_1,
  input      [254:0]  io_inputs_0_payload_state_elements_2,
  input      [254:0]  io_inputs_0_payload_state_elements_3,
  input      [254:0]  io_inputs_0_payload_state_elements_4,
  input      [254:0]  io_inputs_0_payload_state_elements_5,
  input      [254:0]  io_inputs_0_payload_state_elements_6,
  input      [254:0]  io_inputs_0_payload_state_elements_7,
  input      [254:0]  io_inputs_0_payload_state_elements_8,
  input      [254:0]  io_inputs_0_payload_state_elements_9,
  input      [254:0]  io_inputs_0_payload_state_elements_10,
  input      [254:0]  io_inputs_0_payload_state_elements_11,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [6:0]    io_inputs_1_payload_round_index,
  input      [3:0]    io_inputs_1_payload_state_size,
  input      [6:0]    io_inputs_1_payload_state_id,
  input      [254:0]  io_inputs_1_payload_state_elements_0,
  input      [254:0]  io_inputs_1_payload_state_elements_1,
  input      [254:0]  io_inputs_1_payload_state_elements_2,
  input      [254:0]  io_inputs_1_payload_state_elements_3,
  input      [254:0]  io_inputs_1_payload_state_elements_4,
  input      [254:0]  io_inputs_1_payload_state_elements_5,
  input      [254:0]  io_inputs_1_payload_state_elements_6,
  input      [254:0]  io_inputs_1_payload_state_elements_7,
  input      [254:0]  io_inputs_1_payload_state_elements_8,
  input      [254:0]  io_inputs_1_payload_state_elements_9,
  input      [254:0]  io_inputs_1_payload_state_elements_10,
  input      [254:0]  io_inputs_1_payload_state_elements_11,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [6:0]    io_inputs_2_payload_round_index,
  input      [3:0]    io_inputs_2_payload_state_size,
  input      [6:0]    io_inputs_2_payload_state_id,
  input      [254:0]  io_inputs_2_payload_state_elements_0,
  input      [254:0]  io_inputs_2_payload_state_elements_1,
  input      [254:0]  io_inputs_2_payload_state_elements_2,
  input      [254:0]  io_inputs_2_payload_state_elements_3,
  input      [254:0]  io_inputs_2_payload_state_elements_4,
  input      [254:0]  io_inputs_2_payload_state_elements_5,
  input      [254:0]  io_inputs_2_payload_state_elements_6,
  input      [254:0]  io_inputs_2_payload_state_elements_7,
  input      [254:0]  io_inputs_2_payload_state_elements_8,
  input      [254:0]  io_inputs_2_payload_state_elements_9,
  input      [254:0]  io_inputs_2_payload_state_elements_10,
  input      [254:0]  io_inputs_2_payload_state_elements_11,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               clk,
  input               reset
);
  wire       [254:0]  modAdder_1_res_o;
  wire       [254:0]  modAdder_2_res_o;
  wire       [254:0]  modAdder_3_res_o;
  wire       [254:0]  modAdder_4_res_o;
  wire       [254:0]  modAdder_5_res_o;
  wire       [254:0]  modAdder_6_res_o;
  wire       [254:0]  modAdder_7_res_o;
  wire       [254:0]  modAdder_8_res_o;
  wire       [254:0]  modAdder_9_res_o;
  wire       [254:0]  modAdder_10_res_o;
  wire       [254:0]  modAdder_11_res_o;
  wire       [254:0]  modAdder_12_res_o;
  wire       [254:0]  modAdder_13_res_o;
  wire       [254:0]  modAdder_14_res_o;
  wire       [254:0]  modAdder_15_res_o;
  wire       [254:0]  modAdder_16_res_o;
  wire       [254:0]  modAdder_17_res_o;
  wire       [254:0]  modAdder_18_res_o;
  wire       [254:0]  modAdder_19_res_o;
  wire       [254:0]  modAdder_20_res_o;
  wire       [254:0]  modAdder_21_res_o;
  wire       [254:0]  modAdder_22_res_o;
  wire       [254:0]  modAdder_23_res_o;
  wire       [254:0]  modAdder_24_res_o;
  wire       [254:0]  modAdder_25_res_o;
  wire       [254:0]  modAdder_26_res_o;
  wire       [254:0]  modAdder_27_res_o;
  wire       [254:0]  modAdder_28_res_o;
  wire       [254:0]  modAdder_29_res_o;
  wire       [254:0]  modAdder_30_res_o;
  wire       [254:0]  modAdder_31_res_o;
  wire       [254:0]  modAdder_32_res_o;
  wire       [254:0]  modAdder_33_res_o;
  wire       [254:0]  modAdder_34_res_o;
  wire       [254:0]  modAdder_35_res_o;
  wire       [254:0]  modAdder_36_res_o;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l94;
  wire                threadAdders_tempRes_valid;
  reg                 threadAdders_tempRes_ready;
  wire       [6:0]    threadAdders_tempRes_payload_round_index;
  wire       [3:0]    threadAdders_tempRes_payload_state_size;
  wire       [6:0]    threadAdders_tempRes_payload_state_id;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_0;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_1;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_2;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_3;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_4;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_5;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_6;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_7;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_8;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_9;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_10;
  reg        [254:0]  threadAdders_tempRes_payload_state_elements_11;
  wire                _zz_io_inputs_0_ready;
  wire                _zz_io_inputs_0_ready_1;
  wire                threadAdders_tempRes_tempOp1s_valid;
  wire                threadAdders_tempRes_tempOp1s_ready;
  wire       [6:0]    threadAdders_tempRes_tempOp1s_payload_round_index;
  wire       [3:0]    threadAdders_tempRes_tempOp1s_payload_state_size;
  wire       [6:0]    threadAdders_tempRes_tempOp1s_payload_state_id;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_0;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_1;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_2;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_3;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_4;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_5;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_6;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_7;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_8;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_9;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_10;
  wire       [254:0]  threadAdders_tempRes_tempOp1s_payload_state_elements_11;
  reg                 threadAdders_tempRes_rValid;
  reg        [6:0]    threadAdders_tempRes_rData_round_index;
  reg        [3:0]    threadAdders_tempRes_rData_state_size;
  reg        [6:0]    threadAdders_tempRes_rData_state_id;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_0;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_1;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_2;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_3;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_4;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_5;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_6;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_7;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_8;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_9;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_10;
  reg        [254:0]  threadAdders_tempRes_rData_state_elements_11;
  wire                when_Stream_l342;
  wire                threadAdders_tempRes_fire;
  reg        [254:0]  threadAdders_tempOp2s_0;
  reg        [254:0]  threadAdders_tempOp2s_1;
  reg        [254:0]  threadAdders_tempOp2s_2;
  reg        [254:0]  threadAdders_tempOp2s_3;
  reg        [254:0]  threadAdders_tempOp2s_4;
  reg        [254:0]  threadAdders_tempOp2s_5;
  reg        [254:0]  threadAdders_tempOp2s_6;
  reg        [254:0]  threadAdders_tempOp2s_7;
  reg        [254:0]  threadAdders_tempOp2s_8;
  reg        [254:0]  threadAdders_tempOp2s_9;
  reg        [254:0]  threadAdders_tempOp2s_10;
  reg        [254:0]  threadAdders_tempOp2s_11;
  wire                threadAdders_output_valid;
  reg                 threadAdders_output_ready;
  wire       [6:0]    threadAdders_output_payload_round_index;
  wire       [3:0]    threadAdders_output_payload_state_size;
  wire       [6:0]    threadAdders_output_payload_state_id;
  reg        [254:0]  threadAdders_output_payload_state_elements_0;
  reg        [254:0]  threadAdders_output_payload_state_elements_1;
  reg        [254:0]  threadAdders_output_payload_state_elements_2;
  reg        [254:0]  threadAdders_output_payload_state_elements_3;
  reg        [254:0]  threadAdders_output_payload_state_elements_4;
  reg        [254:0]  threadAdders_output_payload_state_elements_5;
  reg        [254:0]  threadAdders_output_payload_state_elements_6;
  reg        [254:0]  threadAdders_output_payload_state_elements_7;
  reg        [254:0]  threadAdders_output_payload_state_elements_8;
  reg        [254:0]  threadAdders_output_payload_state_elements_9;
  reg        [254:0]  threadAdders_output_payload_state_elements_10;
  reg        [254:0]  threadAdders_output_payload_state_elements_11;
  wire                threadAdders_output_input_valid;
  reg                 threadAdders_output_input_ready;
  wire       [6:0]    threadAdders_output_input_payload_round_index;
  wire       [3:0]    threadAdders_output_input_payload_state_size;
  wire       [6:0]    threadAdders_output_input_payload_state_id;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_0;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_1;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_2;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_3;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_4;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_5;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_6;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_7;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_8;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_9;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_10;
  wire       [254:0]  threadAdders_output_input_payload_state_elements_11;
  reg                 threadAdders_output_rValid;
  reg        [6:0]    threadAdders_output_rData_round_index;
  reg        [3:0]    threadAdders_output_rData_state_size;
  reg        [6:0]    threadAdders_output_rData_state_id;
  reg        [254:0]  threadAdders_output_rData_state_elements_0;
  reg        [254:0]  threadAdders_output_rData_state_elements_1;
  reg        [254:0]  threadAdders_output_rData_state_elements_2;
  reg        [254:0]  threadAdders_output_rData_state_elements_3;
  reg        [254:0]  threadAdders_output_rData_state_elements_4;
  reg        [254:0]  threadAdders_output_rData_state_elements_5;
  reg        [254:0]  threadAdders_output_rData_state_elements_6;
  reg        [254:0]  threadAdders_output_rData_state_elements_7;
  reg        [254:0]  threadAdders_output_rData_state_elements_8;
  reg        [254:0]  threadAdders_output_rData_state_elements_9;
  reg        [254:0]  threadAdders_output_rData_state_elements_10;
  reg        [254:0]  threadAdders_output_rData_state_elements_11;
  wire                when_Stream_l342_1;
  reg                 threadAccumulator_output_valid;
  wire                threadAccumulator_output_ready;
  wire       [6:0]    threadAccumulator_output_payload_round_index;
  wire       [3:0]    threadAccumulator_output_payload_state_size;
  wire       [6:0]    threadAccumulator_output_payload_state_id;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_0;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_1;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_2;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_3;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_4;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_5;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_6;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_7;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_8;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_9;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_10;
  wire       [254:0]  threadAccumulator_output_payload_state_elements_11;
  reg        [6:0]    threadAccumulator_tempRes_round_index;
  reg        [3:0]    threadAccumulator_tempRes_state_size;
  reg        [6:0]    threadAccumulator_tempRes_state_id;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_0;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_1;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_2;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_3;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_4;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_5;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_6;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_7;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_8;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_9;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_10;
  reg        [254:0]  threadAccumulator_tempRes_state_elements_11;
  wire       [254:0]  threadAccumulator_modAdderRes_0;
  wire       [254:0]  threadAccumulator_modAdderRes_1;
  wire       [254:0]  threadAccumulator_modAdderRes_2;
  wire       [254:0]  threadAccumulator_modAdderRes_3;
  wire       [254:0]  threadAccumulator_modAdderRes_4;
  wire       [254:0]  threadAccumulator_modAdderRes_5;
  wire       [254:0]  threadAccumulator_modAdderRes_6;
  wire       [254:0]  threadAccumulator_modAdderRes_7;
  wire       [254:0]  threadAccumulator_modAdderRes_8;
  wire       [254:0]  threadAccumulator_modAdderRes_9;
  wire       [254:0]  threadAccumulator_modAdderRes_10;
  wire       [254:0]  threadAccumulator_modAdderRes_11;
  wire                threadAccumulator_fsm_wantExit;
  reg                 threadAccumulator_fsm_wantStart;
  wire                threadAccumulator_fsm_wantKill;
  reg        [3:0]    threadAccumulator_fsm_counter;
  reg        `threadAccumulator_fsm_enumDefinition_binary_sequential_type threadAccumulator_fsm_stateReg;
  reg        `threadAccumulator_fsm_enumDefinition_binary_sequential_type threadAccumulator_fsm_stateNext;
  wire                threadAdders_output_input_fire;
  wire                when_MDSMatrixAdders_l79;
  wire                threadAdders_output_input_fire_1;
  wire                when_MDSMatrixAdders_l94;
  wire                threadAccumulator_output_fire;
  wire                threadAdders_output_input_fire_2;
  wire                when_MDSMatrixAdders_l111;
  wire                when_StateMachine_l214;
  `ifndef SYNTHESIS
  reg [223:0] threadAccumulator_fsm_stateReg_string;
  reg [223:0] threadAccumulator_fsm_stateNext_string;
  `endif


  assign _zz_when_MDSMatrixAdders_l94 = (threadAccumulator_fsm_counter + 4'b0011);
  ModAdder modAdder_1 (
    .op1_i    (io_inputs_0_payload_state_elements_0  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_0  ), //i
    .res_o    (modAdder_1_res_o                      )  //o
  );
  ModAdder modAdder_2 (
    .op1_i    (io_inputs_0_payload_state_elements_1  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_1  ), //i
    .res_o    (modAdder_2_res_o                      )  //o
  );
  ModAdder modAdder_3 (
    .op1_i    (io_inputs_0_payload_state_elements_2  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_2  ), //i
    .res_o    (modAdder_3_res_o                      )  //o
  );
  ModAdder modAdder_4 (
    .op1_i    (io_inputs_0_payload_state_elements_3  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_3  ), //i
    .res_o    (modAdder_4_res_o                      )  //o
  );
  ModAdder modAdder_5 (
    .op1_i    (io_inputs_0_payload_state_elements_4  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_4  ), //i
    .res_o    (modAdder_5_res_o                      )  //o
  );
  ModAdder modAdder_6 (
    .op1_i    (io_inputs_0_payload_state_elements_5  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_5  ), //i
    .res_o    (modAdder_6_res_o                      )  //o
  );
  ModAdder modAdder_7 (
    .op1_i    (io_inputs_0_payload_state_elements_6  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_6  ), //i
    .res_o    (modAdder_7_res_o                      )  //o
  );
  ModAdder modAdder_8 (
    .op1_i    (io_inputs_0_payload_state_elements_7  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_7  ), //i
    .res_o    (modAdder_8_res_o                      )  //o
  );
  ModAdder modAdder_9 (
    .op1_i    (io_inputs_0_payload_state_elements_8  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_8  ), //i
    .res_o    (modAdder_9_res_o                      )  //o
  );
  ModAdder modAdder_10 (
    .op1_i    (io_inputs_0_payload_state_elements_9  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_9  ), //i
    .res_o    (modAdder_10_res_o                     )  //o
  );
  ModAdder modAdder_11 (
    .op1_i    (io_inputs_0_payload_state_elements_10  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_10  ), //i
    .res_o    (modAdder_11_res_o                      )  //o
  );
  ModAdder modAdder_12 (
    .op1_i    (io_inputs_0_payload_state_elements_11  ), //i
    .op2_i    (io_inputs_1_payload_state_elements_11  ), //i
    .res_o    (modAdder_12_res_o                      )  //o
  );
  ModAdder modAdder_13 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_0  ), //i
    .op2_i    (threadAdders_tempOp2s_0                                 ), //i
    .res_o    (modAdder_13_res_o                                       )  //o
  );
  ModAdder modAdder_14 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_1  ), //i
    .op2_i    (threadAdders_tempOp2s_1                                 ), //i
    .res_o    (modAdder_14_res_o                                       )  //o
  );
  ModAdder modAdder_15 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_2  ), //i
    .op2_i    (threadAdders_tempOp2s_2                                 ), //i
    .res_o    (modAdder_15_res_o                                       )  //o
  );
  ModAdder modAdder_16 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_3  ), //i
    .op2_i    (threadAdders_tempOp2s_3                                 ), //i
    .res_o    (modAdder_16_res_o                                       )  //o
  );
  ModAdder modAdder_17 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_4  ), //i
    .op2_i    (threadAdders_tempOp2s_4                                 ), //i
    .res_o    (modAdder_17_res_o                                       )  //o
  );
  ModAdder modAdder_18 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_5  ), //i
    .op2_i    (threadAdders_tempOp2s_5                                 ), //i
    .res_o    (modAdder_18_res_o                                       )  //o
  );
  ModAdder modAdder_19 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_6  ), //i
    .op2_i    (threadAdders_tempOp2s_6                                 ), //i
    .res_o    (modAdder_19_res_o                                       )  //o
  );
  ModAdder modAdder_20 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_7  ), //i
    .op2_i    (threadAdders_tempOp2s_7                                 ), //i
    .res_o    (modAdder_20_res_o                                       )  //o
  );
  ModAdder modAdder_21 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_8  ), //i
    .op2_i    (threadAdders_tempOp2s_8                                 ), //i
    .res_o    (modAdder_21_res_o                                       )  //o
  );
  ModAdder modAdder_22 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_9  ), //i
    .op2_i    (threadAdders_tempOp2s_9                                 ), //i
    .res_o    (modAdder_22_res_o                                       )  //o
  );
  ModAdder modAdder_23 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_10  ), //i
    .op2_i    (threadAdders_tempOp2s_10                                 ), //i
    .res_o    (modAdder_23_res_o                                        )  //o
  );
  ModAdder modAdder_24 (
    .op1_i    (threadAdders_tempRes_tempOp1s_payload_state_elements_11  ), //i
    .op2_i    (threadAdders_tempOp2s_11                                 ), //i
    .res_o    (modAdder_24_res_o                                        )  //o
  );
  ModAdder modAdder_25 (
    .op1_i    (threadAccumulator_tempRes_state_elements_0          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_0  ), //i
    .res_o    (modAdder_25_res_o                                   )  //o
  );
  ModAdder modAdder_26 (
    .op1_i    (threadAccumulator_tempRes_state_elements_1          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_1  ), //i
    .res_o    (modAdder_26_res_o                                   )  //o
  );
  ModAdder modAdder_27 (
    .op1_i    (threadAccumulator_tempRes_state_elements_2          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_2  ), //i
    .res_o    (modAdder_27_res_o                                   )  //o
  );
  ModAdder modAdder_28 (
    .op1_i    (threadAccumulator_tempRes_state_elements_3          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_3  ), //i
    .res_o    (modAdder_28_res_o                                   )  //o
  );
  ModAdder modAdder_29 (
    .op1_i    (threadAccumulator_tempRes_state_elements_4          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_4  ), //i
    .res_o    (modAdder_29_res_o                                   )  //o
  );
  ModAdder modAdder_30 (
    .op1_i    (threadAccumulator_tempRes_state_elements_5          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_5  ), //i
    .res_o    (modAdder_30_res_o                                   )  //o
  );
  ModAdder modAdder_31 (
    .op1_i    (threadAccumulator_tempRes_state_elements_6          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_6  ), //i
    .res_o    (modAdder_31_res_o                                   )  //o
  );
  ModAdder modAdder_32 (
    .op1_i    (threadAccumulator_tempRes_state_elements_7          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_7  ), //i
    .res_o    (modAdder_32_res_o                                   )  //o
  );
  ModAdder modAdder_33 (
    .op1_i    (threadAccumulator_tempRes_state_elements_8          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_8  ), //i
    .res_o    (modAdder_33_res_o                                   )  //o
  );
  ModAdder modAdder_34 (
    .op1_i    (threadAccumulator_tempRes_state_elements_9          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_9  ), //i
    .res_o    (modAdder_34_res_o                                   )  //o
  );
  ModAdder modAdder_35 (
    .op1_i    (threadAccumulator_tempRes_state_elements_10          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_10  ), //i
    .res_o    (modAdder_35_res_o                                    )  //o
  );
  ModAdder modAdder_36 (
    .op1_i    (threadAccumulator_tempRes_state_elements_11          ), //i
    .op2_i    (threadAdders_output_input_payload_state_elements_11  ), //i
    .res_o    (modAdder_36_res_o                                    )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(threadAccumulator_fsm_stateReg)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_BOOT : threadAccumulator_fsm_stateReg_string = "threadAccumulator_fsm_BOOT  ";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : threadAccumulator_fsm_stateReg_string = "threadAccumulator_fsm_IDLE  ";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : threadAccumulator_fsm_stateReg_string = "threadAccumulator_fsm_ADDING";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : threadAccumulator_fsm_stateReg_string = "threadAccumulator_fsm_DONE  ";
      default : threadAccumulator_fsm_stateReg_string = "????????????????????????????";
    endcase
  end
  always @(*) begin
    case(threadAccumulator_fsm_stateNext)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_BOOT : threadAccumulator_fsm_stateNext_string = "threadAccumulator_fsm_BOOT  ";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : threadAccumulator_fsm_stateNext_string = "threadAccumulator_fsm_IDLE  ";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : threadAccumulator_fsm_stateNext_string = "threadAccumulator_fsm_ADDING";
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : threadAccumulator_fsm_stateNext_string = "threadAccumulator_fsm_DONE  ";
      default : threadAccumulator_fsm_stateNext_string = "????????????????????????????";
    endcase
  end
  `endif

  assign _zz_io_inputs_0_ready_1 = (_zz_io_inputs_0_ready && threadAdders_tempRes_ready);
  assign _zz_io_inputs_0_ready = ((io_inputs_0_valid && io_inputs_1_valid) && io_inputs_2_valid);
  assign io_inputs_0_ready = _zz_io_inputs_0_ready_1;
  assign io_inputs_1_ready = _zz_io_inputs_0_ready_1;
  assign io_inputs_2_ready = _zz_io_inputs_0_ready_1;
  assign threadAdders_tempRes_valid = _zz_io_inputs_0_ready;
  assign threadAdders_tempRes_payload_round_index = io_inputs_0_payload_round_index;
  assign threadAdders_tempRes_payload_state_size = io_inputs_0_payload_state_size;
  assign threadAdders_tempRes_payload_state_id = io_inputs_0_payload_state_id;
  always @(*) begin
    threadAdders_tempRes_payload_state_elements_0 = io_inputs_0_payload_state_elements_0;
    threadAdders_tempRes_payload_state_elements_0 = modAdder_1_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_1 = io_inputs_0_payload_state_elements_1;
    threadAdders_tempRes_payload_state_elements_1 = modAdder_2_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_2 = io_inputs_0_payload_state_elements_2;
    threadAdders_tempRes_payload_state_elements_2 = modAdder_3_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_3 = io_inputs_0_payload_state_elements_3;
    threadAdders_tempRes_payload_state_elements_3 = modAdder_4_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_4 = io_inputs_0_payload_state_elements_4;
    threadAdders_tempRes_payload_state_elements_4 = modAdder_5_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_5 = io_inputs_0_payload_state_elements_5;
    threadAdders_tempRes_payload_state_elements_5 = modAdder_6_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_6 = io_inputs_0_payload_state_elements_6;
    threadAdders_tempRes_payload_state_elements_6 = modAdder_7_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_7 = io_inputs_0_payload_state_elements_7;
    threadAdders_tempRes_payload_state_elements_7 = modAdder_8_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_8 = io_inputs_0_payload_state_elements_8;
    threadAdders_tempRes_payload_state_elements_8 = modAdder_9_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_9 = io_inputs_0_payload_state_elements_9;
    threadAdders_tempRes_payload_state_elements_9 = modAdder_10_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_10 = io_inputs_0_payload_state_elements_10;
    threadAdders_tempRes_payload_state_elements_10 = modAdder_11_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_payload_state_elements_11 = io_inputs_0_payload_state_elements_11;
    threadAdders_tempRes_payload_state_elements_11 = modAdder_12_res_o;
  end

  always @(*) begin
    threadAdders_tempRes_ready = threadAdders_tempRes_tempOp1s_ready;
    if(when_Stream_l342) begin
      threadAdders_tempRes_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! threadAdders_tempRes_tempOp1s_valid);
  assign threadAdders_tempRes_tempOp1s_valid = threadAdders_tempRes_rValid;
  assign threadAdders_tempRes_tempOp1s_payload_round_index = threadAdders_tempRes_rData_round_index;
  assign threadAdders_tempRes_tempOp1s_payload_state_size = threadAdders_tempRes_rData_state_size;
  assign threadAdders_tempRes_tempOp1s_payload_state_id = threadAdders_tempRes_rData_state_id;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_0 = threadAdders_tempRes_rData_state_elements_0;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_1 = threadAdders_tempRes_rData_state_elements_1;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_2 = threadAdders_tempRes_rData_state_elements_2;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_3 = threadAdders_tempRes_rData_state_elements_3;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_4 = threadAdders_tempRes_rData_state_elements_4;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_5 = threadAdders_tempRes_rData_state_elements_5;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_6 = threadAdders_tempRes_rData_state_elements_6;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_7 = threadAdders_tempRes_rData_state_elements_7;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_8 = threadAdders_tempRes_rData_state_elements_8;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_9 = threadAdders_tempRes_rData_state_elements_9;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_10 = threadAdders_tempRes_rData_state_elements_10;
  assign threadAdders_tempRes_tempOp1s_payload_state_elements_11 = threadAdders_tempRes_rData_state_elements_11;
  assign threadAdders_tempRes_fire = (threadAdders_tempRes_valid && threadAdders_tempRes_ready);
  assign threadAdders_output_valid = threadAdders_tempRes_tempOp1s_valid;
  assign threadAdders_tempRes_tempOp1s_ready = threadAdders_output_ready;
  assign threadAdders_output_payload_round_index = threadAdders_tempRes_tempOp1s_payload_round_index;
  assign threadAdders_output_payload_state_size = threadAdders_tempRes_tempOp1s_payload_state_size;
  assign threadAdders_output_payload_state_id = threadAdders_tempRes_tempOp1s_payload_state_id;
  always @(*) begin
    threadAdders_output_payload_state_elements_0 = threadAdders_tempRes_tempOp1s_payload_state_elements_0;
    threadAdders_output_payload_state_elements_0 = modAdder_13_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_1 = threadAdders_tempRes_tempOp1s_payload_state_elements_1;
    threadAdders_output_payload_state_elements_1 = modAdder_14_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_2 = threadAdders_tempRes_tempOp1s_payload_state_elements_2;
    threadAdders_output_payload_state_elements_2 = modAdder_15_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_3 = threadAdders_tempRes_tempOp1s_payload_state_elements_3;
    threadAdders_output_payload_state_elements_3 = modAdder_16_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_4 = threadAdders_tempRes_tempOp1s_payload_state_elements_4;
    threadAdders_output_payload_state_elements_4 = modAdder_17_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_5 = threadAdders_tempRes_tempOp1s_payload_state_elements_5;
    threadAdders_output_payload_state_elements_5 = modAdder_18_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_6 = threadAdders_tempRes_tempOp1s_payload_state_elements_6;
    threadAdders_output_payload_state_elements_6 = modAdder_19_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_7 = threadAdders_tempRes_tempOp1s_payload_state_elements_7;
    threadAdders_output_payload_state_elements_7 = modAdder_20_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_8 = threadAdders_tempRes_tempOp1s_payload_state_elements_8;
    threadAdders_output_payload_state_elements_8 = modAdder_21_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_9 = threadAdders_tempRes_tempOp1s_payload_state_elements_9;
    threadAdders_output_payload_state_elements_9 = modAdder_22_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_10 = threadAdders_tempRes_tempOp1s_payload_state_elements_10;
    threadAdders_output_payload_state_elements_10 = modAdder_23_res_o;
  end

  always @(*) begin
    threadAdders_output_payload_state_elements_11 = threadAdders_tempRes_tempOp1s_payload_state_elements_11;
    threadAdders_output_payload_state_elements_11 = modAdder_24_res_o;
  end

  always @(*) begin
    threadAdders_output_ready = threadAdders_output_input_ready;
    if(when_Stream_l342_1) begin
      threadAdders_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! threadAdders_output_input_valid);
  assign threadAdders_output_input_valid = threadAdders_output_rValid;
  assign threadAdders_output_input_payload_round_index = threadAdders_output_rData_round_index;
  assign threadAdders_output_input_payload_state_size = threadAdders_output_rData_state_size;
  assign threadAdders_output_input_payload_state_id = threadAdders_output_rData_state_id;
  assign threadAdders_output_input_payload_state_elements_0 = threadAdders_output_rData_state_elements_0;
  assign threadAdders_output_input_payload_state_elements_1 = threadAdders_output_rData_state_elements_1;
  assign threadAdders_output_input_payload_state_elements_2 = threadAdders_output_rData_state_elements_2;
  assign threadAdders_output_input_payload_state_elements_3 = threadAdders_output_rData_state_elements_3;
  assign threadAdders_output_input_payload_state_elements_4 = threadAdders_output_rData_state_elements_4;
  assign threadAdders_output_input_payload_state_elements_5 = threadAdders_output_rData_state_elements_5;
  assign threadAdders_output_input_payload_state_elements_6 = threadAdders_output_rData_state_elements_6;
  assign threadAdders_output_input_payload_state_elements_7 = threadAdders_output_rData_state_elements_7;
  assign threadAdders_output_input_payload_state_elements_8 = threadAdders_output_rData_state_elements_8;
  assign threadAdders_output_input_payload_state_elements_9 = threadAdders_output_rData_state_elements_9;
  assign threadAdders_output_input_payload_state_elements_10 = threadAdders_output_rData_state_elements_10;
  assign threadAdders_output_input_payload_state_elements_11 = threadAdders_output_rData_state_elements_11;
  assign threadAccumulator_modAdderRes_0 = modAdder_25_res_o;
  assign threadAccumulator_modAdderRes_1 = modAdder_26_res_o;
  assign threadAccumulator_modAdderRes_2 = modAdder_27_res_o;
  assign threadAccumulator_modAdderRes_3 = modAdder_28_res_o;
  assign threadAccumulator_modAdderRes_4 = modAdder_29_res_o;
  assign threadAccumulator_modAdderRes_5 = modAdder_30_res_o;
  assign threadAccumulator_modAdderRes_6 = modAdder_31_res_o;
  assign threadAccumulator_modAdderRes_7 = modAdder_32_res_o;
  assign threadAccumulator_modAdderRes_8 = modAdder_33_res_o;
  assign threadAccumulator_modAdderRes_9 = modAdder_34_res_o;
  assign threadAccumulator_modAdderRes_10 = modAdder_35_res_o;
  assign threadAccumulator_modAdderRes_11 = modAdder_36_res_o;
  assign threadAccumulator_fsm_wantExit = 1'b0;
  always @(*) begin
    threadAccumulator_fsm_wantStart = 1'b0;
    case(threadAccumulator_fsm_stateReg)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : begin
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : begin
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : begin
      end
      default : begin
        threadAccumulator_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign threadAccumulator_fsm_wantKill = 1'b0;
  assign threadAccumulator_output_payload_round_index = threadAccumulator_tempRes_round_index;
  assign threadAccumulator_output_payload_state_size = threadAccumulator_tempRes_state_size;
  assign threadAccumulator_output_payload_state_id = threadAccumulator_tempRes_state_id;
  assign threadAccumulator_output_payload_state_elements_0 = threadAccumulator_tempRes_state_elements_0;
  assign threadAccumulator_output_payload_state_elements_1 = threadAccumulator_tempRes_state_elements_1;
  assign threadAccumulator_output_payload_state_elements_2 = threadAccumulator_tempRes_state_elements_2;
  assign threadAccumulator_output_payload_state_elements_3 = threadAccumulator_tempRes_state_elements_3;
  assign threadAccumulator_output_payload_state_elements_4 = threadAccumulator_tempRes_state_elements_4;
  assign threadAccumulator_output_payload_state_elements_5 = threadAccumulator_tempRes_state_elements_5;
  assign threadAccumulator_output_payload_state_elements_6 = threadAccumulator_tempRes_state_elements_6;
  assign threadAccumulator_output_payload_state_elements_7 = threadAccumulator_tempRes_state_elements_7;
  assign threadAccumulator_output_payload_state_elements_8 = threadAccumulator_tempRes_state_elements_8;
  assign threadAccumulator_output_payload_state_elements_9 = threadAccumulator_tempRes_state_elements_9;
  assign threadAccumulator_output_payload_state_elements_10 = threadAccumulator_tempRes_state_elements_10;
  assign threadAccumulator_output_payload_state_elements_11 = threadAccumulator_tempRes_state_elements_11;
  always @(*) begin
    threadAccumulator_output_valid = 1'b0;
    case(threadAccumulator_fsm_stateReg)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : begin
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : begin
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : begin
        threadAccumulator_output_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    threadAdders_output_input_ready = 1'b0;
    case(threadAccumulator_fsm_stateReg)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : begin
        threadAdders_output_input_ready = 1'b1;
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : begin
        threadAdders_output_input_ready = 1'b1;
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : begin
        if(threadAccumulator_output_fire) begin
          threadAdders_output_input_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign io_output_valid = threadAccumulator_output_valid;
  assign threadAccumulator_output_ready = io_output_ready;
  assign io_output_payload_round_index = threadAccumulator_output_payload_round_index;
  assign io_output_payload_state_size = threadAccumulator_output_payload_state_size;
  assign io_output_payload_state_id = threadAccumulator_output_payload_state_id;
  assign io_output_payload_state_elements_0 = threadAccumulator_output_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = threadAccumulator_output_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = threadAccumulator_output_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = threadAccumulator_output_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = threadAccumulator_output_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = threadAccumulator_output_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = threadAccumulator_output_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = threadAccumulator_output_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = threadAccumulator_output_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = threadAccumulator_output_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = threadAccumulator_output_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = threadAccumulator_output_payload_state_elements_11;
  always @(*) begin
    threadAccumulator_fsm_stateNext = threadAccumulator_fsm_stateReg;
    case(threadAccumulator_fsm_stateReg)
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : begin
        if(threadAdders_output_input_fire) begin
          if(when_MDSMatrixAdders_l79) begin
            threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE;
          end else begin
            threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING;
          end
        end
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : begin
        if(threadAdders_output_input_fire_1) begin
          if(when_MDSMatrixAdders_l94) begin
            threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE;
          end
        end
      end
      `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : begin
        if(threadAccumulator_output_fire) begin
          if(threadAdders_output_input_fire_2) begin
            if(when_MDSMatrixAdders_l111) begin
              threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING;
            end
          end else begin
            threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE;
          end
        end
      end
      default : begin
      end
    endcase
    if(threadAccumulator_fsm_wantStart) begin
      threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE;
    end
    if(threadAccumulator_fsm_wantKill) begin
      threadAccumulator_fsm_stateNext = `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_BOOT;
    end
  end

  assign threadAdders_output_input_fire = (threadAdders_output_input_valid && threadAdders_output_input_ready);
  assign when_MDSMatrixAdders_l79 = (threadAdders_output_input_payload_state_size == 4'b0011);
  assign threadAdders_output_input_fire_1 = (threadAdders_output_input_valid && threadAdders_output_input_ready);
  assign when_MDSMatrixAdders_l94 = (threadAccumulator_tempRes_state_size <= _zz_when_MDSMatrixAdders_l94);
  assign threadAccumulator_output_fire = (threadAccumulator_output_valid && threadAccumulator_output_ready);
  assign threadAdders_output_input_fire_2 = (threadAdders_output_input_valid && threadAdders_output_input_ready);
  assign when_MDSMatrixAdders_l111 = (4'b0011 < threadAdders_output_input_payload_state_size);
  assign when_StateMachine_l214 = ((threadAccumulator_fsm_stateReg == `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING) && (! (threadAccumulator_fsm_stateNext == `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING)));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      threadAdders_tempRes_rValid <= 1'b0;
      threadAdders_tempOp2s_0 <= 255'h0;
      threadAdders_tempOp2s_1 <= 255'h0;
      threadAdders_tempOp2s_2 <= 255'h0;
      threadAdders_tempOp2s_3 <= 255'h0;
      threadAdders_tempOp2s_4 <= 255'h0;
      threadAdders_tempOp2s_5 <= 255'h0;
      threadAdders_tempOp2s_6 <= 255'h0;
      threadAdders_tempOp2s_7 <= 255'h0;
      threadAdders_tempOp2s_8 <= 255'h0;
      threadAdders_tempOp2s_9 <= 255'h0;
      threadAdders_tempOp2s_10 <= 255'h0;
      threadAdders_tempOp2s_11 <= 255'h0;
      threadAdders_output_rValid <= 1'b0;
      threadAccumulator_tempRes_state_size <= 4'b0000;
      threadAccumulator_tempRes_state_elements_0 <= 255'h0;
      threadAccumulator_tempRes_state_elements_1 <= 255'h0;
      threadAccumulator_tempRes_state_elements_2 <= 255'h0;
      threadAccumulator_tempRes_state_elements_3 <= 255'h0;
      threadAccumulator_tempRes_state_elements_4 <= 255'h0;
      threadAccumulator_tempRes_state_elements_5 <= 255'h0;
      threadAccumulator_tempRes_state_elements_6 <= 255'h0;
      threadAccumulator_tempRes_state_elements_7 <= 255'h0;
      threadAccumulator_tempRes_state_elements_8 <= 255'h0;
      threadAccumulator_tempRes_state_elements_9 <= 255'h0;
      threadAccumulator_tempRes_state_elements_10 <= 255'h0;
      threadAccumulator_tempRes_state_elements_11 <= 255'h0;
      threadAccumulator_tempRes_state_id <= 7'h0;
      threadAccumulator_tempRes_round_index <= 7'h0;
      threadAccumulator_fsm_counter <= 4'b0000;
      threadAccumulator_fsm_stateReg <= `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_BOOT;
    end else begin
      if(threadAdders_tempRes_ready) begin
        threadAdders_tempRes_rValid <= threadAdders_tempRes_valid;
      end
      if(threadAdders_tempRes_fire) begin
        threadAdders_tempOp2s_0 <= io_inputs_2_payload_state_elements_0;
        threadAdders_tempOp2s_1 <= io_inputs_2_payload_state_elements_1;
        threadAdders_tempOp2s_2 <= io_inputs_2_payload_state_elements_2;
        threadAdders_tempOp2s_3 <= io_inputs_2_payload_state_elements_3;
        threadAdders_tempOp2s_4 <= io_inputs_2_payload_state_elements_4;
        threadAdders_tempOp2s_5 <= io_inputs_2_payload_state_elements_5;
        threadAdders_tempOp2s_6 <= io_inputs_2_payload_state_elements_6;
        threadAdders_tempOp2s_7 <= io_inputs_2_payload_state_elements_7;
        threadAdders_tempOp2s_8 <= io_inputs_2_payload_state_elements_8;
        threadAdders_tempOp2s_9 <= io_inputs_2_payload_state_elements_9;
        threadAdders_tempOp2s_10 <= io_inputs_2_payload_state_elements_10;
        threadAdders_tempOp2s_11 <= io_inputs_2_payload_state_elements_11;
      end
      if(threadAdders_output_ready) begin
        threadAdders_output_rValid <= threadAdders_output_valid;
      end
      threadAccumulator_fsm_stateReg <= threadAccumulator_fsm_stateNext;
      case(threadAccumulator_fsm_stateReg)
        `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_IDLE : begin
          if(threadAdders_output_input_fire) begin
            threadAccumulator_tempRes_round_index <= threadAdders_output_input_payload_round_index;
            threadAccumulator_tempRes_state_size <= threadAdders_output_input_payload_state_size;
            threadAccumulator_tempRes_state_id <= threadAdders_output_input_payload_state_id;
            threadAccumulator_tempRes_state_elements_0 <= threadAdders_output_input_payload_state_elements_0;
            threadAccumulator_tempRes_state_elements_1 <= threadAdders_output_input_payload_state_elements_1;
            threadAccumulator_tempRes_state_elements_2 <= threadAdders_output_input_payload_state_elements_2;
            threadAccumulator_tempRes_state_elements_3 <= threadAdders_output_input_payload_state_elements_3;
            threadAccumulator_tempRes_state_elements_4 <= threadAdders_output_input_payload_state_elements_4;
            threadAccumulator_tempRes_state_elements_5 <= threadAdders_output_input_payload_state_elements_5;
            threadAccumulator_tempRes_state_elements_6 <= threadAdders_output_input_payload_state_elements_6;
            threadAccumulator_tempRes_state_elements_7 <= threadAdders_output_input_payload_state_elements_7;
            threadAccumulator_tempRes_state_elements_8 <= threadAdders_output_input_payload_state_elements_8;
            threadAccumulator_tempRes_state_elements_9 <= threadAdders_output_input_payload_state_elements_9;
            threadAccumulator_tempRes_state_elements_10 <= threadAdders_output_input_payload_state_elements_10;
            threadAccumulator_tempRes_state_elements_11 <= threadAdders_output_input_payload_state_elements_11;
            if(!when_MDSMatrixAdders_l79) begin
              threadAccumulator_fsm_counter <= (threadAccumulator_fsm_counter + 4'b0011);
            end
          end
        end
        `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_ADDING : begin
          if(threadAdders_output_input_fire_1) begin
            threadAccumulator_tempRes_state_elements_0 <= threadAccumulator_modAdderRes_0;
            threadAccumulator_tempRes_state_elements_1 <= threadAccumulator_modAdderRes_1;
            threadAccumulator_tempRes_state_elements_2 <= threadAccumulator_modAdderRes_2;
            threadAccumulator_tempRes_state_elements_3 <= threadAccumulator_modAdderRes_3;
            threadAccumulator_tempRes_state_elements_4 <= threadAccumulator_modAdderRes_4;
            threadAccumulator_tempRes_state_elements_5 <= threadAccumulator_modAdderRes_5;
            threadAccumulator_tempRes_state_elements_6 <= threadAccumulator_modAdderRes_6;
            threadAccumulator_tempRes_state_elements_7 <= threadAccumulator_modAdderRes_7;
            threadAccumulator_tempRes_state_elements_8 <= threadAccumulator_modAdderRes_8;
            threadAccumulator_tempRes_state_elements_9 <= threadAccumulator_modAdderRes_9;
            threadAccumulator_tempRes_state_elements_10 <= threadAccumulator_modAdderRes_10;
            threadAccumulator_tempRes_state_elements_11 <= threadAccumulator_modAdderRes_11;
            if(!when_MDSMatrixAdders_l94) begin
              threadAccumulator_fsm_counter <= (threadAccumulator_fsm_counter + 4'b0011);
            end
          end
        end
        `threadAccumulator_fsm_enumDefinition_binary_sequential_threadAccumulator_fsm_DONE : begin
          if(threadAccumulator_output_fire) begin
            if(threadAdders_output_input_fire_2) begin
              threadAccumulator_tempRes_round_index <= threadAdders_output_input_payload_round_index;
              threadAccumulator_tempRes_state_size <= threadAdders_output_input_payload_state_size;
              threadAccumulator_tempRes_state_id <= threadAdders_output_input_payload_state_id;
              threadAccumulator_tempRes_state_elements_0 <= threadAdders_output_input_payload_state_elements_0;
              threadAccumulator_tempRes_state_elements_1 <= threadAdders_output_input_payload_state_elements_1;
              threadAccumulator_tempRes_state_elements_2 <= threadAdders_output_input_payload_state_elements_2;
              threadAccumulator_tempRes_state_elements_3 <= threadAdders_output_input_payload_state_elements_3;
              threadAccumulator_tempRes_state_elements_4 <= threadAdders_output_input_payload_state_elements_4;
              threadAccumulator_tempRes_state_elements_5 <= threadAdders_output_input_payload_state_elements_5;
              threadAccumulator_tempRes_state_elements_6 <= threadAdders_output_input_payload_state_elements_6;
              threadAccumulator_tempRes_state_elements_7 <= threadAdders_output_input_payload_state_elements_7;
              threadAccumulator_tempRes_state_elements_8 <= threadAdders_output_input_payload_state_elements_8;
              threadAccumulator_tempRes_state_elements_9 <= threadAdders_output_input_payload_state_elements_9;
              threadAccumulator_tempRes_state_elements_10 <= threadAdders_output_input_payload_state_elements_10;
              threadAccumulator_tempRes_state_elements_11 <= threadAdders_output_input_payload_state_elements_11;
              if(when_MDSMatrixAdders_l111) begin
                threadAccumulator_fsm_counter <= (threadAccumulator_fsm_counter + 4'b0011);
              end
            end
          end
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l214) begin
        threadAccumulator_fsm_counter <= 4'b0000;
      end
    end
  end

  always @(posedge clk) begin
    if(threadAdders_tempRes_ready) begin
      threadAdders_tempRes_rData_round_index <= threadAdders_tempRes_payload_round_index;
      threadAdders_tempRes_rData_state_size <= threadAdders_tempRes_payload_state_size;
      threadAdders_tempRes_rData_state_id <= threadAdders_tempRes_payload_state_id;
      threadAdders_tempRes_rData_state_elements_0 <= threadAdders_tempRes_payload_state_elements_0;
      threadAdders_tempRes_rData_state_elements_1 <= threadAdders_tempRes_payload_state_elements_1;
      threadAdders_tempRes_rData_state_elements_2 <= threadAdders_tempRes_payload_state_elements_2;
      threadAdders_tempRes_rData_state_elements_3 <= threadAdders_tempRes_payload_state_elements_3;
      threadAdders_tempRes_rData_state_elements_4 <= threadAdders_tempRes_payload_state_elements_4;
      threadAdders_tempRes_rData_state_elements_5 <= threadAdders_tempRes_payload_state_elements_5;
      threadAdders_tempRes_rData_state_elements_6 <= threadAdders_tempRes_payload_state_elements_6;
      threadAdders_tempRes_rData_state_elements_7 <= threadAdders_tempRes_payload_state_elements_7;
      threadAdders_tempRes_rData_state_elements_8 <= threadAdders_tempRes_payload_state_elements_8;
      threadAdders_tempRes_rData_state_elements_9 <= threadAdders_tempRes_payload_state_elements_9;
      threadAdders_tempRes_rData_state_elements_10 <= threadAdders_tempRes_payload_state_elements_10;
      threadAdders_tempRes_rData_state_elements_11 <= threadAdders_tempRes_payload_state_elements_11;
    end
    if(threadAdders_output_ready) begin
      threadAdders_output_rData_round_index <= threadAdders_output_payload_round_index;
      threadAdders_output_rData_state_size <= threadAdders_output_payload_state_size;
      threadAdders_output_rData_state_id <= threadAdders_output_payload_state_id;
      threadAdders_output_rData_state_elements_0 <= threadAdders_output_payload_state_elements_0;
      threadAdders_output_rData_state_elements_1 <= threadAdders_output_payload_state_elements_1;
      threadAdders_output_rData_state_elements_2 <= threadAdders_output_payload_state_elements_2;
      threadAdders_output_rData_state_elements_3 <= threadAdders_output_payload_state_elements_3;
      threadAdders_output_rData_state_elements_4 <= threadAdders_output_payload_state_elements_4;
      threadAdders_output_rData_state_elements_5 <= threadAdders_output_payload_state_elements_5;
      threadAdders_output_rData_state_elements_6 <= threadAdders_output_payload_state_elements_6;
      threadAdders_output_rData_state_elements_7 <= threadAdders_output_payload_state_elements_7;
      threadAdders_output_rData_state_elements_8 <= threadAdders_output_payload_state_elements_8;
      threadAdders_output_rData_state_elements_9 <= threadAdders_output_payload_state_elements_9;
      threadAdders_output_rData_state_elements_10 <= threadAdders_output_payload_state_elements_10;
      threadAdders_output_rData_state_elements_11 <= threadAdders_output_payload_state_elements_11;
    end
  end


endmodule

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

module AXI4StreamReceiver (
  input               io_input_valid,
  output reg          io_input_ready,
  input               io_input_last,
  input      [254:0]  io_input_payload,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_round_index,
  output     [3:0]    io_outputs_0_payload_state_index,
  output     [3:0]    io_outputs_0_payload_state_size,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [254:0]  io_outputs_0_payload_state_element,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_round_index,
  output     [3:0]    io_outputs_1_payload_state_index,
  output     [3:0]    io_outputs_1_payload_state_size,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [254:0]  io_outputs_1_payload_state_element,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [6:0]    io_outputs_2_payload_round_index,
  output     [3:0]    io_outputs_2_payload_state_index,
  output     [3:0]    io_outputs_2_payload_state_size,
  output     [6:0]    io_outputs_2_payload_state_id,
  output     [254:0]  io_outputs_2_payload_state_element,
  input               clk,
  input               reset
);
  wire                DataBuffer_buffer2_buffer3_buffer3_fork_io_input_ready;
  wire                DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_valid;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_round_index;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_size;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_id;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_2;
  wire                DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_valid;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_round_index;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_size;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_id;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_2;
  wire                DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_valid;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_round_index;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_size;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_id;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_2;
  reg        [6:0]    DataController_idCounter;
  reg        [3:0]    DataController_lengthCounter;
  reg        [254:0]  DataController_state_elements_0;
  reg        [254:0]  DataController_state_elements_1;
  reg        [254:0]  DataController_state_elements_2;
  reg        [3:0]    DataController_state_indexes_0;
  reg        [3:0]    DataController_state_indexes_1;
  reg        [3:0]    DataController_state_indexes_2;
  reg                 DataController_output_valid;
  reg                 DataController_output_ready;
  wire       [6:0]    DataController_output_payload_round_index;
  wire       [3:0]    DataController_output_payload_state_size;
  wire       [6:0]    DataController_output_payload_state_id;
  wire       [3:0]    DataController_output_payload_state_indexes_0;
  wire       [3:0]    DataController_output_payload_state_indexes_1;
  wire       [3:0]    DataController_output_payload_state_indexes_2;
  wire       [254:0]  DataController_output_payload_state_elements_0;
  wire       [254:0]  DataController_output_payload_state_elements_1;
  wire       [254:0]  DataController_output_payload_state_elements_2;
  reg        `ReceiverState_binary_sequential_type DataController_receiverState;
  wire                when_AXI4StreamInterface_l52;
  wire                when_AXI4StreamInterface_l63;
  wire                when_AXI4StreamInterface_l79;
  wire                DataController_output_fire;
  wire                when_AXI4StreamInterface_l99;
  wire                when_AXI4StreamInterface_l114;
  wire                DataController_output_fire_1;
  wire                when_AXI4StreamInterface_l131;
  wire                DataBuffer_continue;
  wire                DataController_output_buffer0_valid;
  wire                DataController_output_buffer0_ready;
  wire       [6:0]    DataController_output_buffer0_payload_round_index;
  wire       [3:0]    DataController_output_buffer0_payload_state_size;
  wire       [6:0]    DataController_output_buffer0_payload_state_id;
  wire       [3:0]    DataController_output_buffer0_payload_state_indexes_0;
  wire       [3:0]    DataController_output_buffer0_payload_state_indexes_1;
  wire       [3:0]    DataController_output_buffer0_payload_state_indexes_2;
  wire       [254:0]  DataController_output_buffer0_payload_state_elements_0;
  wire       [254:0]  DataController_output_buffer0_payload_state_elements_1;
  wire       [254:0]  DataController_output_buffer0_payload_state_elements_2;
  reg                 DataController_output_rValid;
  reg        [6:0]    DataController_output_rData_round_index;
  reg        [3:0]    DataController_output_rData_state_size;
  reg        [6:0]    DataController_output_rData_state_id;
  reg        [3:0]    DataController_output_rData_state_indexes_0;
  reg        [3:0]    DataController_output_rData_state_indexes_1;
  reg        [3:0]    DataController_output_rData_state_indexes_2;
  reg        [254:0]  DataController_output_rData_state_elements_0;
  reg        [254:0]  DataController_output_rData_state_elements_1;
  reg        [254:0]  DataController_output_rData_state_elements_2;
  wire                when_Stream_l342;
  wire                DataBuffer_buffer0_buffer1_valid;
  reg                 DataBuffer_buffer0_buffer1_ready;
  wire       [6:0]    DataBuffer_buffer0_buffer1_payload_round_index;
  reg        [3:0]    DataBuffer_buffer0_buffer1_payload_state_size;
  wire       [6:0]    DataBuffer_buffer0_buffer1_payload_state_id;
  wire       [3:0]    DataBuffer_buffer0_buffer1_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer0_buffer1_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer0_buffer1_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer0_buffer1_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer0_buffer1_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer0_buffer1_payload_state_elements_2;
  wire                _zz_DataController_output_buffer0_ready;
  wire                when_AXI4StreamInterface_l155;
  wire                when_AXI4StreamInterface_l156;
  wire                DataBuffer_buffer0_buffer1_buffer1_valid;
  wire                DataBuffer_buffer0_buffer1_buffer1_ready;
  wire       [6:0]    DataBuffer_buffer0_buffer1_buffer1_payload_round_index;
  wire       [3:0]    DataBuffer_buffer0_buffer1_buffer1_payload_state_size;
  wire       [6:0]    DataBuffer_buffer0_buffer1_buffer1_payload_state_id;
  wire       [3:0]    DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_2;
  reg                 DataBuffer_buffer0_buffer1_rValid;
  reg        [6:0]    DataBuffer_buffer0_buffer1_rData_round_index;
  reg        [3:0]    DataBuffer_buffer0_buffer1_rData_state_size;
  reg        [6:0]    DataBuffer_buffer0_buffer1_rData_state_id;
  reg        [3:0]    DataBuffer_buffer0_buffer1_rData_state_indexes_0;
  reg        [3:0]    DataBuffer_buffer0_buffer1_rData_state_indexes_1;
  reg        [3:0]    DataBuffer_buffer0_buffer1_rData_state_indexes_2;
  reg        [254:0]  DataBuffer_buffer0_buffer1_rData_state_elements_0;
  reg        [254:0]  DataBuffer_buffer0_buffer1_rData_state_elements_1;
  reg        [254:0]  DataBuffer_buffer0_buffer1_rData_state_elements_2;
  wire                when_Stream_l342_1;
  wire                DataBuffer_buffer1_buffer2_valid;
  reg                 DataBuffer_buffer1_buffer2_ready;
  wire       [6:0]    DataBuffer_buffer1_buffer2_payload_round_index;
  reg        [3:0]    DataBuffer_buffer1_buffer2_payload_state_size;
  wire       [6:0]    DataBuffer_buffer1_buffer2_payload_state_id;
  wire       [3:0]    DataBuffer_buffer1_buffer2_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer1_buffer2_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer1_buffer2_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer1_buffer2_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer1_buffer2_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer1_buffer2_payload_state_elements_2;
  wire                _zz_DataBuffer_buffer0_buffer1_buffer1_ready;
  wire                when_AXI4StreamInterface_l167;
  wire                when_AXI4StreamInterface_l168;
  wire                DataBuffer_buffer1_buffer2_buffer2_valid;
  wire                DataBuffer_buffer1_buffer2_buffer2_ready;
  wire       [6:0]    DataBuffer_buffer1_buffer2_buffer2_payload_round_index;
  wire       [3:0]    DataBuffer_buffer1_buffer2_buffer2_payload_state_size;
  wire       [6:0]    DataBuffer_buffer1_buffer2_buffer2_payload_state_id;
  wire       [3:0]    DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_2;
  reg                 DataBuffer_buffer1_buffer2_rValid;
  reg        [6:0]    DataBuffer_buffer1_buffer2_rData_round_index;
  reg        [3:0]    DataBuffer_buffer1_buffer2_rData_state_size;
  reg        [6:0]    DataBuffer_buffer1_buffer2_rData_state_id;
  reg        [3:0]    DataBuffer_buffer1_buffer2_rData_state_indexes_0;
  reg        [3:0]    DataBuffer_buffer1_buffer2_rData_state_indexes_1;
  reg        [3:0]    DataBuffer_buffer1_buffer2_rData_state_indexes_2;
  reg        [254:0]  DataBuffer_buffer1_buffer2_rData_state_elements_0;
  reg        [254:0]  DataBuffer_buffer1_buffer2_rData_state_elements_1;
  reg        [254:0]  DataBuffer_buffer1_buffer2_rData_state_elements_2;
  wire                when_Stream_l342_2;
  wire                DataBuffer_buffer2_buffer3_valid;
  reg                 DataBuffer_buffer2_buffer3_ready;
  wire       [6:0]    DataBuffer_buffer2_buffer3_payload_round_index;
  reg        [3:0]    DataBuffer_buffer2_buffer3_payload_state_size;
  wire       [6:0]    DataBuffer_buffer2_buffer3_payload_state_id;
  wire       [3:0]    DataBuffer_buffer2_buffer3_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer2_buffer3_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer2_buffer3_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer2_buffer3_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer2_buffer3_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer2_buffer3_payload_state_elements_2;
  wire                _zz_DataBuffer_buffer1_buffer2_buffer2_ready;
  wire                when_AXI4StreamInterface_l179;
  wire                when_AXI4StreamInterface_l180;
  wire                DataBuffer_buffer2_buffer3_buffer3_valid;
  wire                DataBuffer_buffer2_buffer3_buffer3_ready;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_payload_round_index;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_payload_state_size;
  wire       [6:0]    DataBuffer_buffer2_buffer3_buffer3_payload_state_id;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_0;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_1;
  wire       [3:0]    DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_2;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_0;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_1;
  wire       [254:0]  DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_2;
  reg                 DataBuffer_buffer2_buffer3_rValid;
  reg        [6:0]    DataBuffer_buffer2_buffer3_rData_round_index;
  reg        [3:0]    DataBuffer_buffer2_buffer3_rData_state_size;
  reg        [6:0]    DataBuffer_buffer2_buffer3_rData_state_id;
  reg        [3:0]    DataBuffer_buffer2_buffer3_rData_state_indexes_0;
  reg        [3:0]    DataBuffer_buffer2_buffer3_rData_state_indexes_1;
  reg        [3:0]    DataBuffer_buffer2_buffer3_rData_state_indexes_2;
  reg        [254:0]  DataBuffer_buffer2_buffer3_rData_state_elements_0;
  reg        [254:0]  DataBuffer_buffer2_buffer3_rData_state_elements_1;
  reg        [254:0]  DataBuffer_buffer2_buffer3_rData_state_elements_2;
  wire                when_Stream_l342_3;
  `ifndef SYNTHESIS
  reg [79:0] DataController_receiverState_string;
  `endif


  StreamFork_9 DataBuffer_buffer2_buffer3_buffer3_fork (
    .io_input_valid                           (DataBuffer_buffer2_buffer3_buffer3_valid                                       ), //i
    .io_input_ready                           (DataBuffer_buffer2_buffer3_buffer3_fork_io_input_ready                         ), //o
    .io_input_payload_round_index             (DataBuffer_buffer2_buffer3_buffer3_payload_round_index                         ), //i
    .io_input_payload_state_size              (DataBuffer_buffer2_buffer3_buffer3_payload_state_size                          ), //i
    .io_input_payload_state_id                (DataBuffer_buffer2_buffer3_buffer3_payload_state_id                            ), //i
    .io_input_payload_state_indexes_0         (DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_0                     ), //i
    .io_input_payload_state_indexes_1         (DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_1                     ), //i
    .io_input_payload_state_indexes_2         (DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_2                     ), //i
    .io_input_payload_state_elements_0        (DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_0                    ), //i
    .io_input_payload_state_elements_1        (DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_1                    ), //i
    .io_input_payload_state_elements_2        (DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_2                    ), //i
    .io_outputs_0_valid                       (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_valid                     ), //o
    .io_outputs_0_ready                       (io_outputs_0_ready                                                             ), //i
    .io_outputs_0_payload_round_index         (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_round_index       ), //o
    .io_outputs_0_payload_state_size          (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_size        ), //o
    .io_outputs_0_payload_state_id            (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_id          ), //o
    .io_outputs_0_payload_state_indexes_0     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_0   ), //o
    .io_outputs_0_payload_state_indexes_1     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_1   ), //o
    .io_outputs_0_payload_state_indexes_2     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_2   ), //o
    .io_outputs_0_payload_state_elements_0    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_0  ), //o
    .io_outputs_0_payload_state_elements_1    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_1  ), //o
    .io_outputs_0_payload_state_elements_2    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_2  ), //o
    .io_outputs_1_valid                       (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_valid                     ), //o
    .io_outputs_1_ready                       (io_outputs_1_ready                                                             ), //i
    .io_outputs_1_payload_round_index         (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_round_index       ), //o
    .io_outputs_1_payload_state_size          (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_size        ), //o
    .io_outputs_1_payload_state_id            (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_id          ), //o
    .io_outputs_1_payload_state_indexes_0     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_0   ), //o
    .io_outputs_1_payload_state_indexes_1     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_1   ), //o
    .io_outputs_1_payload_state_indexes_2     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_2   ), //o
    .io_outputs_1_payload_state_elements_0    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_0  ), //o
    .io_outputs_1_payload_state_elements_1    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_1  ), //o
    .io_outputs_1_payload_state_elements_2    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_2  ), //o
    .io_outputs_2_valid                       (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_valid                     ), //o
    .io_outputs_2_ready                       (io_outputs_2_ready                                                             ), //i
    .io_outputs_2_payload_round_index         (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_round_index       ), //o
    .io_outputs_2_payload_state_size          (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_size        ), //o
    .io_outputs_2_payload_state_id            (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_id          ), //o
    .io_outputs_2_payload_state_indexes_0     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_0   ), //o
    .io_outputs_2_payload_state_indexes_1     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_1   ), //o
    .io_outputs_2_payload_state_indexes_2     (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_2   ), //o
    .io_outputs_2_payload_state_elements_0    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_0  ), //o
    .io_outputs_2_payload_state_elements_1    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_1  ), //o
    .io_outputs_2_payload_state_elements_2    (DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_2  )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(DataController_receiverState)
      `ReceiverState_binary_sequential_IDLE : DataController_receiverState_string = "IDLE      ";
      `ReceiverState_binary_sequential_ELEMENT0 : DataController_receiverState_string = "ELEMENT0  ";
      `ReceiverState_binary_sequential_ELEMENT1 : DataController_receiverState_string = "ELEMENT1  ";
      `ReceiverState_binary_sequential_BLOCK_1 : DataController_receiverState_string = "BLOCK_1   ";
      `ReceiverState_binary_sequential_BLOCK_IDLE : DataController_receiverState_string = "BLOCK_IDLE";
      `ReceiverState_binary_sequential_DONE : DataController_receiverState_string = "DONE      ";
      default : DataController_receiverState_string = "??????????";
    endcase
  end
  `endif

  assign DataController_output_payload_round_index = 7'h0;
  assign DataController_output_payload_state_size = DataController_lengthCounter;
  assign DataController_output_payload_state_id = DataController_idCounter;
  assign DataController_output_payload_state_indexes_0 = DataController_state_indexes_0;
  assign DataController_output_payload_state_indexes_1 = DataController_state_indexes_1;
  assign DataController_output_payload_state_indexes_2 = DataController_state_indexes_2;
  assign DataController_output_payload_state_elements_0 = DataController_state_elements_0;
  assign DataController_output_payload_state_elements_1 = DataController_state_elements_1;
  assign DataController_output_payload_state_elements_2 = DataController_state_elements_2;
  always @(*) begin
    DataController_output_valid = 1'b0;
    case(DataController_receiverState)
      `ReceiverState_binary_sequential_IDLE : begin
      end
      `ReceiverState_binary_sequential_ELEMENT0 : begin
      end
      `ReceiverState_binary_sequential_ELEMENT1 : begin
      end
      `ReceiverState_binary_sequential_BLOCK_1 : begin
        DataController_output_valid = 1'b1;
      end
      `ReceiverState_binary_sequential_BLOCK_IDLE : begin
      end
      default : begin
        DataController_output_valid = 1'b1;
      end
    endcase
  end

  always @(*) begin
    io_input_ready = 1'b0;
    case(DataController_receiverState)
      `ReceiverState_binary_sequential_IDLE : begin
        io_input_ready = 1'b1;
      end
      `ReceiverState_binary_sequential_ELEMENT0 : begin
        io_input_ready = 1'b1;
      end
      `ReceiverState_binary_sequential_ELEMENT1 : begin
        io_input_ready = 1'b1;
      end
      `ReceiverState_binary_sequential_BLOCK_1 : begin
        if(DataController_output_fire) begin
          io_input_ready = 1'b1;
        end
      end
      `ReceiverState_binary_sequential_BLOCK_IDLE : begin
        io_input_ready = 1'b1;
      end
      default : begin
        if(DataController_output_fire_1) begin
          io_input_ready = 1'b1;
        end
      end
    endcase
  end

  assign when_AXI4StreamInterface_l52 = (io_input_valid && io_input_ready);
  assign when_AXI4StreamInterface_l63 = (io_input_valid && io_input_ready);
  assign when_AXI4StreamInterface_l79 = (io_input_valid && io_input_ready);
  assign DataController_output_fire = (DataController_output_valid && DataController_output_ready);
  assign when_AXI4StreamInterface_l99 = (io_input_valid && io_input_ready);
  assign when_AXI4StreamInterface_l114 = (io_input_valid && io_input_ready);
  assign DataController_output_fire_1 = (DataController_output_valid && DataController_output_ready);
  assign when_AXI4StreamInterface_l131 = (io_input_valid && io_input_ready);
  assign DataBuffer_continue = (((DataController_receiverState == `ReceiverState_binary_sequential_DONE) || (DataController_receiverState == `ReceiverState_binary_sequential_BLOCK_1)) || (DataController_receiverState == `ReceiverState_binary_sequential_IDLE));
  always @(*) begin
    DataController_output_ready = DataController_output_buffer0_ready;
    if(when_Stream_l342) begin
      DataController_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! DataController_output_buffer0_valid);
  assign DataController_output_buffer0_valid = DataController_output_rValid;
  assign DataController_output_buffer0_payload_round_index = DataController_output_rData_round_index;
  assign DataController_output_buffer0_payload_state_size = DataController_output_rData_state_size;
  assign DataController_output_buffer0_payload_state_id = DataController_output_rData_state_id;
  assign DataController_output_buffer0_payload_state_indexes_0 = DataController_output_rData_state_indexes_0;
  assign DataController_output_buffer0_payload_state_indexes_1 = DataController_output_rData_state_indexes_1;
  assign DataController_output_buffer0_payload_state_indexes_2 = DataController_output_rData_state_indexes_2;
  assign DataController_output_buffer0_payload_state_elements_0 = DataController_output_rData_state_elements_0;
  assign DataController_output_buffer0_payload_state_elements_1 = DataController_output_rData_state_elements_1;
  assign DataController_output_buffer0_payload_state_elements_2 = DataController_output_rData_state_elements_2;
  assign _zz_DataController_output_buffer0_ready = (DataBuffer_continue || (DataController_output_buffer0_payload_state_id != DataController_idCounter));
  assign DataController_output_buffer0_ready = (DataBuffer_buffer0_buffer1_ready && _zz_DataController_output_buffer0_ready);
  assign DataBuffer_buffer0_buffer1_valid = (DataController_output_buffer0_valid && _zz_DataController_output_buffer0_ready);
  assign DataBuffer_buffer0_buffer1_payload_round_index = DataController_output_buffer0_payload_round_index;
  always @(*) begin
    DataBuffer_buffer0_buffer1_payload_state_size = DataController_output_buffer0_payload_state_size;
    DataBuffer_buffer0_buffer1_payload_state_size = DataController_output_buffer0_payload_state_size;
    if(when_AXI4StreamInterface_l155) begin
      if(when_AXI4StreamInterface_l156) begin
        DataBuffer_buffer0_buffer1_payload_state_size = DataController_lengthCounter;
      end
    end
  end

  assign DataBuffer_buffer0_buffer1_payload_state_id = DataController_output_buffer0_payload_state_id;
  assign DataBuffer_buffer0_buffer1_payload_state_indexes_0 = DataController_output_buffer0_payload_state_indexes_0;
  assign DataBuffer_buffer0_buffer1_payload_state_indexes_1 = DataController_output_buffer0_payload_state_indexes_1;
  assign DataBuffer_buffer0_buffer1_payload_state_indexes_2 = DataController_output_buffer0_payload_state_indexes_2;
  assign DataBuffer_buffer0_buffer1_payload_state_elements_0 = DataController_output_buffer0_payload_state_elements_0;
  assign DataBuffer_buffer0_buffer1_payload_state_elements_1 = DataController_output_buffer0_payload_state_elements_1;
  assign DataBuffer_buffer0_buffer1_payload_state_elements_2 = DataController_output_buffer0_payload_state_elements_2;
  assign when_AXI4StreamInterface_l155 = (DataController_receiverState == `ReceiverState_binary_sequential_DONE);
  assign when_AXI4StreamInterface_l156 = (4'b0011 < DataController_lengthCounter);
  always @(*) begin
    DataBuffer_buffer0_buffer1_ready = DataBuffer_buffer0_buffer1_buffer1_ready;
    if(when_Stream_l342_1) begin
      DataBuffer_buffer0_buffer1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! DataBuffer_buffer0_buffer1_buffer1_valid);
  assign DataBuffer_buffer0_buffer1_buffer1_valid = DataBuffer_buffer0_buffer1_rValid;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_round_index = DataBuffer_buffer0_buffer1_rData_round_index;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_size = DataBuffer_buffer0_buffer1_rData_state_size;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_id = DataBuffer_buffer0_buffer1_rData_state_id;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_0 = DataBuffer_buffer0_buffer1_rData_state_indexes_0;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_1 = DataBuffer_buffer0_buffer1_rData_state_indexes_1;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_2 = DataBuffer_buffer0_buffer1_rData_state_indexes_2;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_0 = DataBuffer_buffer0_buffer1_rData_state_elements_0;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_1 = DataBuffer_buffer0_buffer1_rData_state_elements_1;
  assign DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_2 = DataBuffer_buffer0_buffer1_rData_state_elements_2;
  assign _zz_DataBuffer_buffer0_buffer1_buffer1_ready = (DataBuffer_continue || (DataBuffer_buffer0_buffer1_buffer1_payload_state_id != DataController_idCounter));
  assign DataBuffer_buffer0_buffer1_buffer1_ready = (DataBuffer_buffer1_buffer2_ready && _zz_DataBuffer_buffer0_buffer1_buffer1_ready);
  assign DataBuffer_buffer1_buffer2_valid = (DataBuffer_buffer0_buffer1_buffer1_valid && _zz_DataBuffer_buffer0_buffer1_buffer1_ready);
  assign DataBuffer_buffer1_buffer2_payload_round_index = DataBuffer_buffer0_buffer1_buffer1_payload_round_index;
  always @(*) begin
    DataBuffer_buffer1_buffer2_payload_state_size = DataBuffer_buffer0_buffer1_buffer1_payload_state_size;
    DataBuffer_buffer1_buffer2_payload_state_size = DataBuffer_buffer0_buffer1_buffer1_payload_state_size;
    if(when_AXI4StreamInterface_l167) begin
      if(when_AXI4StreamInterface_l168) begin
        DataBuffer_buffer1_buffer2_payload_state_size = DataController_lengthCounter;
      end
    end
  end

  assign DataBuffer_buffer1_buffer2_payload_state_id = DataBuffer_buffer0_buffer1_buffer1_payload_state_id;
  assign DataBuffer_buffer1_buffer2_payload_state_indexes_0 = DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_0;
  assign DataBuffer_buffer1_buffer2_payload_state_indexes_1 = DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_1;
  assign DataBuffer_buffer1_buffer2_payload_state_indexes_2 = DataBuffer_buffer0_buffer1_buffer1_payload_state_indexes_2;
  assign DataBuffer_buffer1_buffer2_payload_state_elements_0 = DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_0;
  assign DataBuffer_buffer1_buffer2_payload_state_elements_1 = DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_1;
  assign DataBuffer_buffer1_buffer2_payload_state_elements_2 = DataBuffer_buffer0_buffer1_buffer1_payload_state_elements_2;
  assign when_AXI4StreamInterface_l167 = (DataController_receiverState == `ReceiverState_binary_sequential_DONE);
  assign when_AXI4StreamInterface_l168 = (4'b0110 < DataController_lengthCounter);
  always @(*) begin
    DataBuffer_buffer1_buffer2_ready = DataBuffer_buffer1_buffer2_buffer2_ready;
    if(when_Stream_l342_2) begin
      DataBuffer_buffer1_buffer2_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! DataBuffer_buffer1_buffer2_buffer2_valid);
  assign DataBuffer_buffer1_buffer2_buffer2_valid = DataBuffer_buffer1_buffer2_rValid;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_round_index = DataBuffer_buffer1_buffer2_rData_round_index;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_size = DataBuffer_buffer1_buffer2_rData_state_size;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_id = DataBuffer_buffer1_buffer2_rData_state_id;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_0 = DataBuffer_buffer1_buffer2_rData_state_indexes_0;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_1 = DataBuffer_buffer1_buffer2_rData_state_indexes_1;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_2 = DataBuffer_buffer1_buffer2_rData_state_indexes_2;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_0 = DataBuffer_buffer1_buffer2_rData_state_elements_0;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_1 = DataBuffer_buffer1_buffer2_rData_state_elements_1;
  assign DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_2 = DataBuffer_buffer1_buffer2_rData_state_elements_2;
  assign _zz_DataBuffer_buffer1_buffer2_buffer2_ready = (DataBuffer_continue || (DataBuffer_buffer1_buffer2_buffer2_payload_state_id != DataController_idCounter));
  assign DataBuffer_buffer1_buffer2_buffer2_ready = (DataBuffer_buffer2_buffer3_ready && _zz_DataBuffer_buffer1_buffer2_buffer2_ready);
  assign DataBuffer_buffer2_buffer3_valid = (DataBuffer_buffer1_buffer2_buffer2_valid && _zz_DataBuffer_buffer1_buffer2_buffer2_ready);
  assign DataBuffer_buffer2_buffer3_payload_round_index = DataBuffer_buffer1_buffer2_buffer2_payload_round_index;
  always @(*) begin
    DataBuffer_buffer2_buffer3_payload_state_size = DataBuffer_buffer1_buffer2_buffer2_payload_state_size;
    DataBuffer_buffer2_buffer3_payload_state_size = DataBuffer_buffer1_buffer2_buffer2_payload_state_size;
    if(when_AXI4StreamInterface_l179) begin
      if(when_AXI4StreamInterface_l180) begin
        DataBuffer_buffer2_buffer3_payload_state_size = DataController_lengthCounter;
      end
    end
  end

  assign DataBuffer_buffer2_buffer3_payload_state_id = DataBuffer_buffer1_buffer2_buffer2_payload_state_id;
  assign DataBuffer_buffer2_buffer3_payload_state_indexes_0 = DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_0;
  assign DataBuffer_buffer2_buffer3_payload_state_indexes_1 = DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_1;
  assign DataBuffer_buffer2_buffer3_payload_state_indexes_2 = DataBuffer_buffer1_buffer2_buffer2_payload_state_indexes_2;
  assign DataBuffer_buffer2_buffer3_payload_state_elements_0 = DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_0;
  assign DataBuffer_buffer2_buffer3_payload_state_elements_1 = DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_1;
  assign DataBuffer_buffer2_buffer3_payload_state_elements_2 = DataBuffer_buffer1_buffer2_buffer2_payload_state_elements_2;
  assign when_AXI4StreamInterface_l179 = (DataController_receiverState == `ReceiverState_binary_sequential_DONE);
  assign when_AXI4StreamInterface_l180 = (4'b1001 < DataController_lengthCounter);
  always @(*) begin
    DataBuffer_buffer2_buffer3_ready = DataBuffer_buffer2_buffer3_buffer3_ready;
    if(when_Stream_l342_3) begin
      DataBuffer_buffer2_buffer3_ready = 1'b1;
    end
  end

  assign when_Stream_l342_3 = (! DataBuffer_buffer2_buffer3_buffer3_valid);
  assign DataBuffer_buffer2_buffer3_buffer3_valid = DataBuffer_buffer2_buffer3_rValid;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_round_index = DataBuffer_buffer2_buffer3_rData_round_index;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_size = DataBuffer_buffer2_buffer3_rData_state_size;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_id = DataBuffer_buffer2_buffer3_rData_state_id;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_0 = DataBuffer_buffer2_buffer3_rData_state_indexes_0;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_1 = DataBuffer_buffer2_buffer3_rData_state_indexes_1;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_indexes_2 = DataBuffer_buffer2_buffer3_rData_state_indexes_2;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_0 = DataBuffer_buffer2_buffer3_rData_state_elements_0;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_1 = DataBuffer_buffer2_buffer3_rData_state_elements_1;
  assign DataBuffer_buffer2_buffer3_buffer3_payload_state_elements_2 = DataBuffer_buffer2_buffer3_rData_state_elements_2;
  assign DataBuffer_buffer2_buffer3_buffer3_ready = DataBuffer_buffer2_buffer3_buffer3_fork_io_input_ready;
  assign io_outputs_0_valid = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_valid;
  assign io_outputs_0_payload_round_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_round_index;
  assign io_outputs_0_payload_state_size = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_size;
  assign io_outputs_0_payload_state_id = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_id;
  assign io_outputs_0_payload_state_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_indexes_0;
  assign io_outputs_0_payload_state_element = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_0_payload_state_elements_0;
  assign io_outputs_1_valid = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_valid;
  assign io_outputs_1_payload_round_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_round_index;
  assign io_outputs_1_payload_state_size = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_size;
  assign io_outputs_1_payload_state_id = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_id;
  assign io_outputs_1_payload_state_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_indexes_1;
  assign io_outputs_1_payload_state_element = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_1_payload_state_elements_1;
  assign io_outputs_2_valid = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_valid;
  assign io_outputs_2_payload_round_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_round_index;
  assign io_outputs_2_payload_state_size = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_size;
  assign io_outputs_2_payload_state_id = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_id;
  assign io_outputs_2_payload_state_index = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_indexes_2;
  assign io_outputs_2_payload_state_element = DataBuffer_buffer2_buffer3_buffer3_fork_io_outputs_2_payload_state_elements_2;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      DataController_idCounter <= 7'h0;
      DataController_lengthCounter <= 4'b0000;
      DataController_state_elements_0 <= 255'h0;
      DataController_state_elements_1 <= 255'h0;
      DataController_state_elements_2 <= 255'h0;
      DataController_state_indexes_0 <= 4'b0000;
      DataController_state_indexes_1 <= 4'b0000;
      DataController_state_indexes_2 <= 4'b0000;
      DataController_receiverState <= `ReceiverState_binary_sequential_IDLE;
      DataController_output_rValid <= 1'b0;
      DataBuffer_buffer0_buffer1_rValid <= 1'b0;
      DataBuffer_buffer1_buffer2_rValid <= 1'b0;
      DataBuffer_buffer2_buffer3_rValid <= 1'b0;
    end else begin
      case(DataController_receiverState)
        `ReceiverState_binary_sequential_IDLE : begin
          if(when_AXI4StreamInterface_l52) begin
            DataController_state_indexes_0 <= DataController_lengthCounter;
            DataController_state_elements_0 <= io_input_payload;
            DataController_lengthCounter <= (DataController_lengthCounter + 4'b0001);
            DataController_receiverState <= `ReceiverState_binary_sequential_ELEMENT0;
          end
        end
        `ReceiverState_binary_sequential_ELEMENT0 : begin
          if(when_AXI4StreamInterface_l63) begin
            DataController_state_indexes_1 <= DataController_lengthCounter;
            DataController_state_elements_1 <= io_input_payload;
            DataController_lengthCounter <= (DataController_lengthCounter + 4'b0001);
            if(io_input_last) begin
              DataController_state_indexes_2 <= (DataController_lengthCounter + 4'b0001);
              DataController_receiverState <= `ReceiverState_binary_sequential_DONE;
            end else begin
              DataController_receiverState <= `ReceiverState_binary_sequential_ELEMENT1;
            end
          end
        end
        `ReceiverState_binary_sequential_ELEMENT1 : begin
          if(when_AXI4StreamInterface_l79) begin
            DataController_state_indexes_2 <= DataController_lengthCounter;
            DataController_state_elements_2 <= io_input_payload;
            DataController_lengthCounter <= (DataController_lengthCounter + 4'b0001);
            if(io_input_last) begin
              DataController_receiverState <= `ReceiverState_binary_sequential_DONE;
            end else begin
              DataController_receiverState <= `ReceiverState_binary_sequential_BLOCK_1;
            end
          end
        end
        `ReceiverState_binary_sequential_BLOCK_1 : begin
          if(DataController_output_fire) begin
            DataController_state_indexes_0 <= 4'b0000;
            DataController_state_indexes_1 <= 4'b0000;
            DataController_state_indexes_2 <= 4'b0000;
            DataController_state_elements_0 <= 255'h0;
            DataController_state_elements_1 <= 255'h0;
            DataController_state_elements_2 <= 255'h0;
            if(when_AXI4StreamInterface_l99) begin
              DataController_state_indexes_0 <= DataController_lengthCounter;
              DataController_state_elements_0 <= io_input_payload;
              DataController_lengthCounter <= (DataController_lengthCounter + 4'b0001);
              DataController_receiverState <= `ReceiverState_binary_sequential_ELEMENT0;
            end else begin
              DataController_receiverState <= `ReceiverState_binary_sequential_BLOCK_IDLE;
            end
          end
        end
        `ReceiverState_binary_sequential_BLOCK_IDLE : begin
          if(when_AXI4StreamInterface_l114) begin
            DataController_state_indexes_0 <= DataController_lengthCounter;
            DataController_state_elements_0 <= io_input_payload;
            DataController_lengthCounter <= (DataController_lengthCounter + 4'b0001);
            DataController_receiverState <= `ReceiverState_binary_sequential_ELEMENT0;
          end
        end
        default : begin
          if(DataController_output_fire_1) begin
            DataController_lengthCounter <= 4'b0000;
            DataController_idCounter <= (DataController_idCounter + 7'h01);
            DataController_state_indexes_0 <= 4'b0000;
            DataController_state_indexes_1 <= 4'b0000;
            DataController_state_indexes_2 <= 4'b0000;
            DataController_state_elements_0 <= 255'h0;
            DataController_state_elements_1 <= 255'h0;
            DataController_state_elements_2 <= 255'h0;
            if(when_AXI4StreamInterface_l131) begin
              DataController_state_elements_0 <= io_input_payload;
              DataController_lengthCounter <= 4'b0001;
              DataController_receiverState <= `ReceiverState_binary_sequential_ELEMENT0;
            end else begin
              DataController_receiverState <= `ReceiverState_binary_sequential_IDLE;
            end
          end
        end
      endcase
      if(DataController_output_ready) begin
        DataController_output_rValid <= DataController_output_valid;
      end
      if(DataBuffer_buffer0_buffer1_ready) begin
        DataBuffer_buffer0_buffer1_rValid <= DataBuffer_buffer0_buffer1_valid;
      end
      if(DataBuffer_buffer1_buffer2_ready) begin
        DataBuffer_buffer1_buffer2_rValid <= DataBuffer_buffer1_buffer2_valid;
      end
      if(DataBuffer_buffer2_buffer3_ready) begin
        DataBuffer_buffer2_buffer3_rValid <= DataBuffer_buffer2_buffer3_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(DataController_output_ready) begin
      DataController_output_rData_round_index <= DataController_output_payload_round_index;
      DataController_output_rData_state_size <= DataController_output_payload_state_size;
      DataController_output_rData_state_id <= DataController_output_payload_state_id;
      DataController_output_rData_state_indexes_0 <= DataController_output_payload_state_indexes_0;
      DataController_output_rData_state_indexes_1 <= DataController_output_payload_state_indexes_1;
      DataController_output_rData_state_indexes_2 <= DataController_output_payload_state_indexes_2;
      DataController_output_rData_state_elements_0 <= DataController_output_payload_state_elements_0;
      DataController_output_rData_state_elements_1 <= DataController_output_payload_state_elements_1;
      DataController_output_rData_state_elements_2 <= DataController_output_payload_state_elements_2;
    end
    if(DataBuffer_buffer0_buffer1_ready) begin
      DataBuffer_buffer0_buffer1_rData_round_index <= DataBuffer_buffer0_buffer1_payload_round_index;
      DataBuffer_buffer0_buffer1_rData_state_size <= DataBuffer_buffer0_buffer1_payload_state_size;
      DataBuffer_buffer0_buffer1_rData_state_id <= DataBuffer_buffer0_buffer1_payload_state_id;
      DataBuffer_buffer0_buffer1_rData_state_indexes_0 <= DataBuffer_buffer0_buffer1_payload_state_indexes_0;
      DataBuffer_buffer0_buffer1_rData_state_indexes_1 <= DataBuffer_buffer0_buffer1_payload_state_indexes_1;
      DataBuffer_buffer0_buffer1_rData_state_indexes_2 <= DataBuffer_buffer0_buffer1_payload_state_indexes_2;
      DataBuffer_buffer0_buffer1_rData_state_elements_0 <= DataBuffer_buffer0_buffer1_payload_state_elements_0;
      DataBuffer_buffer0_buffer1_rData_state_elements_1 <= DataBuffer_buffer0_buffer1_payload_state_elements_1;
      DataBuffer_buffer0_buffer1_rData_state_elements_2 <= DataBuffer_buffer0_buffer1_payload_state_elements_2;
    end
    if(DataBuffer_buffer1_buffer2_ready) begin
      DataBuffer_buffer1_buffer2_rData_round_index <= DataBuffer_buffer1_buffer2_payload_round_index;
      DataBuffer_buffer1_buffer2_rData_state_size <= DataBuffer_buffer1_buffer2_payload_state_size;
      DataBuffer_buffer1_buffer2_rData_state_id <= DataBuffer_buffer1_buffer2_payload_state_id;
      DataBuffer_buffer1_buffer2_rData_state_indexes_0 <= DataBuffer_buffer1_buffer2_payload_state_indexes_0;
      DataBuffer_buffer1_buffer2_rData_state_indexes_1 <= DataBuffer_buffer1_buffer2_payload_state_indexes_1;
      DataBuffer_buffer1_buffer2_rData_state_indexes_2 <= DataBuffer_buffer1_buffer2_payload_state_indexes_2;
      DataBuffer_buffer1_buffer2_rData_state_elements_0 <= DataBuffer_buffer1_buffer2_payload_state_elements_0;
      DataBuffer_buffer1_buffer2_rData_state_elements_1 <= DataBuffer_buffer1_buffer2_payload_state_elements_1;
      DataBuffer_buffer1_buffer2_rData_state_elements_2 <= DataBuffer_buffer1_buffer2_payload_state_elements_2;
    end
    if(DataBuffer_buffer2_buffer3_ready) begin
      DataBuffer_buffer2_buffer3_rData_round_index <= DataBuffer_buffer2_buffer3_payload_round_index;
      DataBuffer_buffer2_buffer3_rData_state_size <= DataBuffer_buffer2_buffer3_payload_state_size;
      DataBuffer_buffer2_buffer3_rData_state_id <= DataBuffer_buffer2_buffer3_payload_state_id;
      DataBuffer_buffer2_buffer3_rData_state_indexes_0 <= DataBuffer_buffer2_buffer3_payload_state_indexes_0;
      DataBuffer_buffer2_buffer3_rData_state_indexes_1 <= DataBuffer_buffer2_buffer3_payload_state_indexes_1;
      DataBuffer_buffer2_buffer3_rData_state_indexes_2 <= DataBuffer_buffer2_buffer3_payload_state_indexes_2;
      DataBuffer_buffer2_buffer3_rData_state_elements_0 <= DataBuffer_buffer2_buffer3_payload_state_elements_0;
      DataBuffer_buffer2_buffer3_rData_state_elements_1 <= DataBuffer_buffer2_buffer3_payload_state_elements_1;
      DataBuffer_buffer2_buffer3_rData_state_elements_2 <= DataBuffer_buffer2_buffer3_payload_state_elements_2;
    end
  end


endmodule

module StreamMux_6 (
  input      [2:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [6:0]    io_inputs_0_payload_state_id,
  input      [254:0]  io_inputs_0_payload_state_element,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [6:0]    io_inputs_1_payload_state_id,
  input      [254:0]  io_inputs_1_payload_state_element,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [6:0]    io_inputs_2_payload_state_id,
  input      [254:0]  io_inputs_2_payload_state_element,
  input               io_inputs_3_valid,
  output              io_inputs_3_ready,
  input      [6:0]    io_inputs_3_payload_state_id,
  input      [254:0]  io_inputs_3_payload_state_element,
  input               io_inputs_4_valid,
  output              io_inputs_4_ready,
  input      [6:0]    io_inputs_4_payload_state_id,
  input      [254:0]  io_inputs_4_payload_state_element,
  input               io_inputs_5_valid,
  output              io_inputs_5_ready,
  input      [6:0]    io_inputs_5_payload_state_id,
  input      [254:0]  io_inputs_5_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_element
);
  reg                 _zz_io_output_valid;
  reg        [6:0]    _zz_io_output_payload_state_id;
  reg        [254:0]  _zz_io_output_payload_state_element;

  always @(*) begin
    case(io_select)
      3'b000 : begin
        _zz_io_output_valid = io_inputs_0_valid;
        _zz_io_output_payload_state_id = io_inputs_0_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_0_payload_state_element;
      end
      3'b001 : begin
        _zz_io_output_valid = io_inputs_1_valid;
        _zz_io_output_payload_state_id = io_inputs_1_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_1_payload_state_element;
      end
      3'b010 : begin
        _zz_io_output_valid = io_inputs_2_valid;
        _zz_io_output_payload_state_id = io_inputs_2_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_2_payload_state_element;
      end
      3'b011 : begin
        _zz_io_output_valid = io_inputs_3_valid;
        _zz_io_output_payload_state_id = io_inputs_3_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_3_payload_state_element;
      end
      3'b100 : begin
        _zz_io_output_valid = io_inputs_4_valid;
        _zz_io_output_payload_state_id = io_inputs_4_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_4_payload_state_element;
      end
      default : begin
        _zz_io_output_valid = io_inputs_5_valid;
        _zz_io_output_payload_state_id = io_inputs_5_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_5_payload_state_element;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 3'b000) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 3'b001) && io_output_ready);
  assign io_inputs_2_ready = ((io_select == 3'b010) && io_output_ready);
  assign io_inputs_3_ready = ((io_select == 3'b011) && io_output_ready);
  assign io_inputs_4_ready = ((io_select == 3'b100) && io_output_ready);
  assign io_inputs_5_ready = ((io_select == 3'b101) && io_output_ready);
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_state_id = _zz_io_output_payload_state_id;
  assign io_output_payload_state_element = _zz_io_output_payload_state_element;

endmodule

module StreamDemux_6 (
  input      [2:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [254:0]  io_outputs_0_payload_state_element,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [254:0]  io_outputs_1_payload_state_element,
  output reg          io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [6:0]    io_outputs_2_payload_state_id,
  output     [254:0]  io_outputs_2_payload_state_element,
  output reg          io_outputs_3_valid,
  input               io_outputs_3_ready,
  output     [6:0]    io_outputs_3_payload_state_id,
  output     [254:0]  io_outputs_3_payload_state_element,
  output reg          io_outputs_4_valid,
  input               io_outputs_4_ready,
  output     [6:0]    io_outputs_4_payload_state_id,
  output     [254:0]  io_outputs_4_payload_state_element,
  output reg          io_outputs_5_valid,
  input               io_outputs_5_ready,
  output     [6:0]    io_outputs_5_payload_state_id,
  output     [254:0]  io_outputs_5_payload_state_element
);
  wire                when_Stream_l745;
  wire                when_Stream_l745_1;
  wire                when_Stream_l745_2;
  wire                when_Stream_l745_3;
  wire                when_Stream_l745_4;
  wire                when_Stream_l745_5;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l745) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l745_1) begin
      io_input_ready = io_outputs_1_ready;
    end
    if(!when_Stream_l745_2) begin
      io_input_ready = io_outputs_2_ready;
    end
    if(!when_Stream_l745_3) begin
      io_input_ready = io_outputs_3_ready;
    end
    if(!when_Stream_l745_4) begin
      io_input_ready = io_outputs_4_ready;
    end
    if(!when_Stream_l745_5) begin
      io_input_ready = io_outputs_5_ready;
    end
  end

  assign io_outputs_0_payload_state_id = io_input_payload_state_id;
  assign io_outputs_0_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745 = (3'b000 != io_select);
  always @(*) begin
    if(when_Stream_l745) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_state_id = io_input_payload_state_id;
  assign io_outputs_1_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_1 = (3'b001 != io_select);
  always @(*) begin
    if(when_Stream_l745_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end

  assign io_outputs_2_payload_state_id = io_input_payload_state_id;
  assign io_outputs_2_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_2 = (3'b010 != io_select);
  always @(*) begin
    if(when_Stream_l745_2) begin
      io_outputs_2_valid = 1'b0;
    end else begin
      io_outputs_2_valid = io_input_valid;
    end
  end

  assign io_outputs_3_payload_state_id = io_input_payload_state_id;
  assign io_outputs_3_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_3 = (3'b011 != io_select);
  always @(*) begin
    if(when_Stream_l745_3) begin
      io_outputs_3_valid = 1'b0;
    end else begin
      io_outputs_3_valid = io_input_valid;
    end
  end

  assign io_outputs_4_payload_state_id = io_input_payload_state_id;
  assign io_outputs_4_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_4 = (3'b100 != io_select);
  always @(*) begin
    if(when_Stream_l745_4) begin
      io_outputs_4_valid = 1'b0;
    end else begin
      io_outputs_4_valid = io_input_valid;
    end
  end

  assign io_outputs_5_payload_state_id = io_input_payload_state_id;
  assign io_outputs_5_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_5 = (3'b101 != io_select);
  always @(*) begin
    if(when_Stream_l745_5) begin
      io_outputs_5_valid = 1'b0;
    end else begin
      io_outputs_5_valid = io_input_valid;
    end
  end


endmodule

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

//StreamArbiter replaced by StreamArbiter

module StreamArbiter (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [6:0]    io_inputs_0_payload_round_index,
  input      [3:0]    io_inputs_0_payload_state_index,
  input      [3:0]    io_inputs_0_payload_state_size,
  input      [6:0]    io_inputs_0_payload_state_id,
  input      [254:0]  io_inputs_0_payload_state_element,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [6:0]    io_inputs_1_payload_round_index,
  input      [3:0]    io_inputs_1_payload_state_index,
  input      [3:0]    io_inputs_1_payload_state_size,
  input      [6:0]    io_inputs_1_payload_state_id,
  input      [254:0]  io_inputs_1_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_element,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               reset
);
  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_round_index = (maskRouted_0 ? io_inputs_0_payload_round_index : io_inputs_1_payload_round_index);
  assign io_output_payload_state_index = (maskRouted_0 ? io_inputs_0_payload_state_index : io_inputs_1_payload_state_index);
  assign io_output_payload_state_size = (maskRouted_0 ? io_inputs_0_payload_state_size : io_inputs_1_payload_state_size);
  assign io_output_payload_state_id = (maskRouted_0 ? io_inputs_0_payload_state_id : io_inputs_1_payload_state_id);
  assign io_output_payload_state_element = (maskRouted_0 ? io_inputs_0_payload_state_element : io_inputs_1_payload_state_element);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

//StreamMux_1 replaced by StreamMux_1

//StreamFifoLowLatency_1 replaced by StreamFifoLowLatency_1

//StreamDemux replaced by StreamDemux

//StreamFork_10 replaced by StreamFork_10

module MDSMatrixMultiplier_8 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_32 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_33 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_34 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_35 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier_7 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_28 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_29 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_30 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_31 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier_6 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_24 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_25 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_26 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_27 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

//StreamMux replaced by StreamMux

//StreamFifoLowLatency replaced by StreamFifoLowLatency

//StreamDemux replaced by StreamDemux

//StreamFork_10 replaced by StreamFork_10

//SBox5 replaced by SBox5

//SBox5 replaced by SBox5

//SBox5 replaced by SBox5

module RoundConstants_11 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  wire       [254:0]  _zz_constants_roms_9_port0;
  wire       [254:0]  _zz_constants_roms_10_port0;
  wire       [254:0]  _zz_constants_roms_11_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_9 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_10 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_11 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_9.bin",constants_roms_9);
  end
  assign _zz_constants_roms_9_port0 = constants_roms_9[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_10.bin",constants_roms_10);
  end
  assign _zz_constants_roms_10_port0 = constants_roms_10[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t12_constants_roms_11.bin",constants_roms_11);
  end
  assign _zz_constants_roms_11_port0 = constants_roms_11[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      4'b1000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
      4'b1001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_9_port0;
      end
      4'b1010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_10_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_11_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_10 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t9_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_9 (
  output     [254:0]  io_read_ports_0_data,
  input      [2:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:63];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t5_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t5_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t5_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t5_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t5_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      3'b000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      3'b001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      3'b010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      3'b011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_8 (
  output     [254:0]  io_read_ports_0_data,
  input      [1:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:62];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t3_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t3_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_AddRoundConstantStage_roundConstants_t3_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      2'b00 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      2'b01 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

//StreamMux_1 replaced by StreamMux_1

//StreamFifoLowLatency_1 replaced by StreamFifoLowLatency_1

//StreamDemux replaced by StreamDemux

//StreamFork_10 replaced by StreamFork_10

module MDSMatrixMultiplier_5 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_20 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_21 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_22 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_23 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier_4 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_16 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_17 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_18 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_19 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier_3 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_12 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_13 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_14 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_15 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

//StreamMux replaced by StreamMux

//StreamFifoLowLatency replaced by StreamFifoLowLatency

//StreamDemux replaced by StreamDemux

//StreamFork_10 replaced by StreamFork_10

//SBox5 replaced by SBox5

//SBox5 replaced by SBox5

//SBox5 replaced by SBox5

module RoundConstants_7 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  wire       [254:0]  _zz_constants_roms_9_port0;
  wire       [254:0]  _zz_constants_roms_10_port0;
  wire       [254:0]  _zz_constants_roms_11_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_9 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_10 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_11 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_9.bin",constants_roms_9);
  end
  assign _zz_constants_roms_9_port0 = constants_roms_9[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_10.bin",constants_roms_10);
  end
  assign _zz_constants_roms_10_port0 = constants_roms_10[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t12_constants_roms_11.bin",constants_roms_11);
  end
  assign _zz_constants_roms_11_port0 = constants_roms_11[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      4'b1000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
      4'b1001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_9_port0;
      end
      4'b1010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_10_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_11_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_6 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t9_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_5 (
  output     [254:0]  io_read_ports_0_data,
  input      [2:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:63];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t5_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t5_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t5_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t5_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t5_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      3'b000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      3'b001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      3'b010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      3'b011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_4 (
  output     [254:0]  io_read_ports_0_data,
  input      [1:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:62];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t3_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t3_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_AddRoundConstantStage_roundConstants_t3_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      2'b00 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      2'b01 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module StreamMux_1 (
  input      [1:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [6:0]    io_inputs_0_payload_round_index,
  input      [3:0]    io_inputs_0_payload_state_size,
  input      [6:0]    io_inputs_0_payload_state_id,
  input      [254:0]  io_inputs_0_payload_state_elements_0,
  input      [254:0]  io_inputs_0_payload_state_elements_1,
  input      [254:0]  io_inputs_0_payload_state_elements_2,
  input      [254:0]  io_inputs_0_payload_state_elements_3,
  input      [254:0]  io_inputs_0_payload_state_elements_4,
  input      [254:0]  io_inputs_0_payload_state_elements_5,
  input      [254:0]  io_inputs_0_payload_state_elements_6,
  input      [254:0]  io_inputs_0_payload_state_elements_7,
  input      [254:0]  io_inputs_0_payload_state_elements_8,
  input      [254:0]  io_inputs_0_payload_state_elements_9,
  input      [254:0]  io_inputs_0_payload_state_elements_10,
  input      [254:0]  io_inputs_0_payload_state_elements_11,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [6:0]    io_inputs_1_payload_round_index,
  input      [3:0]    io_inputs_1_payload_state_size,
  input      [6:0]    io_inputs_1_payload_state_id,
  input      [254:0]  io_inputs_1_payload_state_elements_0,
  input      [254:0]  io_inputs_1_payload_state_elements_1,
  input      [254:0]  io_inputs_1_payload_state_elements_2,
  input      [254:0]  io_inputs_1_payload_state_elements_3,
  input      [254:0]  io_inputs_1_payload_state_elements_4,
  input      [254:0]  io_inputs_1_payload_state_elements_5,
  input      [254:0]  io_inputs_1_payload_state_elements_6,
  input      [254:0]  io_inputs_1_payload_state_elements_7,
  input      [254:0]  io_inputs_1_payload_state_elements_8,
  input      [254:0]  io_inputs_1_payload_state_elements_9,
  input      [254:0]  io_inputs_1_payload_state_elements_10,
  input      [254:0]  io_inputs_1_payload_state_elements_11,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [6:0]    io_inputs_2_payload_round_index,
  input      [3:0]    io_inputs_2_payload_state_size,
  input      [6:0]    io_inputs_2_payload_state_id,
  input      [254:0]  io_inputs_2_payload_state_elements_0,
  input      [254:0]  io_inputs_2_payload_state_elements_1,
  input      [254:0]  io_inputs_2_payload_state_elements_2,
  input      [254:0]  io_inputs_2_payload_state_elements_3,
  input      [254:0]  io_inputs_2_payload_state_elements_4,
  input      [254:0]  io_inputs_2_payload_state_elements_5,
  input      [254:0]  io_inputs_2_payload_state_elements_6,
  input      [254:0]  io_inputs_2_payload_state_elements_7,
  input      [254:0]  io_inputs_2_payload_state_elements_8,
  input      [254:0]  io_inputs_2_payload_state_elements_9,
  input      [254:0]  io_inputs_2_payload_state_elements_10,
  input      [254:0]  io_inputs_2_payload_state_elements_11,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11
);
  reg                 _zz_io_output_valid;
  reg        [6:0]    _zz_io_output_payload_round_index;
  reg        [3:0]    _zz_io_output_payload_state_size;
  reg        [6:0]    _zz_io_output_payload_state_id;
  reg        [254:0]  _zz_io_output_payload_state_elements_0;
  reg        [254:0]  _zz_io_output_payload_state_elements_1;
  reg        [254:0]  _zz_io_output_payload_state_elements_2;
  reg        [254:0]  _zz_io_output_payload_state_elements_3;
  reg        [254:0]  _zz_io_output_payload_state_elements_4;
  reg        [254:0]  _zz_io_output_payload_state_elements_5;
  reg        [254:0]  _zz_io_output_payload_state_elements_6;
  reg        [254:0]  _zz_io_output_payload_state_elements_7;
  reg        [254:0]  _zz_io_output_payload_state_elements_8;
  reg        [254:0]  _zz_io_output_payload_state_elements_9;
  reg        [254:0]  _zz_io_output_payload_state_elements_10;
  reg        [254:0]  _zz_io_output_payload_state_elements_11;

  always @(*) begin
    case(io_select)
      2'b00 : begin
        _zz_io_output_valid = io_inputs_0_valid;
        _zz_io_output_payload_round_index = io_inputs_0_payload_round_index;
        _zz_io_output_payload_state_size = io_inputs_0_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_0_payload_state_id;
        _zz_io_output_payload_state_elements_0 = io_inputs_0_payload_state_elements_0;
        _zz_io_output_payload_state_elements_1 = io_inputs_0_payload_state_elements_1;
        _zz_io_output_payload_state_elements_2 = io_inputs_0_payload_state_elements_2;
        _zz_io_output_payload_state_elements_3 = io_inputs_0_payload_state_elements_3;
        _zz_io_output_payload_state_elements_4 = io_inputs_0_payload_state_elements_4;
        _zz_io_output_payload_state_elements_5 = io_inputs_0_payload_state_elements_5;
        _zz_io_output_payload_state_elements_6 = io_inputs_0_payload_state_elements_6;
        _zz_io_output_payload_state_elements_7 = io_inputs_0_payload_state_elements_7;
        _zz_io_output_payload_state_elements_8 = io_inputs_0_payload_state_elements_8;
        _zz_io_output_payload_state_elements_9 = io_inputs_0_payload_state_elements_9;
        _zz_io_output_payload_state_elements_10 = io_inputs_0_payload_state_elements_10;
        _zz_io_output_payload_state_elements_11 = io_inputs_0_payload_state_elements_11;
      end
      2'b01 : begin
        _zz_io_output_valid = io_inputs_1_valid;
        _zz_io_output_payload_round_index = io_inputs_1_payload_round_index;
        _zz_io_output_payload_state_size = io_inputs_1_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_1_payload_state_id;
        _zz_io_output_payload_state_elements_0 = io_inputs_1_payload_state_elements_0;
        _zz_io_output_payload_state_elements_1 = io_inputs_1_payload_state_elements_1;
        _zz_io_output_payload_state_elements_2 = io_inputs_1_payload_state_elements_2;
        _zz_io_output_payload_state_elements_3 = io_inputs_1_payload_state_elements_3;
        _zz_io_output_payload_state_elements_4 = io_inputs_1_payload_state_elements_4;
        _zz_io_output_payload_state_elements_5 = io_inputs_1_payload_state_elements_5;
        _zz_io_output_payload_state_elements_6 = io_inputs_1_payload_state_elements_6;
        _zz_io_output_payload_state_elements_7 = io_inputs_1_payload_state_elements_7;
        _zz_io_output_payload_state_elements_8 = io_inputs_1_payload_state_elements_8;
        _zz_io_output_payload_state_elements_9 = io_inputs_1_payload_state_elements_9;
        _zz_io_output_payload_state_elements_10 = io_inputs_1_payload_state_elements_10;
        _zz_io_output_payload_state_elements_11 = io_inputs_1_payload_state_elements_11;
      end
      default : begin
        _zz_io_output_valid = io_inputs_2_valid;
        _zz_io_output_payload_round_index = io_inputs_2_payload_round_index;
        _zz_io_output_payload_state_size = io_inputs_2_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_2_payload_state_id;
        _zz_io_output_payload_state_elements_0 = io_inputs_2_payload_state_elements_0;
        _zz_io_output_payload_state_elements_1 = io_inputs_2_payload_state_elements_1;
        _zz_io_output_payload_state_elements_2 = io_inputs_2_payload_state_elements_2;
        _zz_io_output_payload_state_elements_3 = io_inputs_2_payload_state_elements_3;
        _zz_io_output_payload_state_elements_4 = io_inputs_2_payload_state_elements_4;
        _zz_io_output_payload_state_elements_5 = io_inputs_2_payload_state_elements_5;
        _zz_io_output_payload_state_elements_6 = io_inputs_2_payload_state_elements_6;
        _zz_io_output_payload_state_elements_7 = io_inputs_2_payload_state_elements_7;
        _zz_io_output_payload_state_elements_8 = io_inputs_2_payload_state_elements_8;
        _zz_io_output_payload_state_elements_9 = io_inputs_2_payload_state_elements_9;
        _zz_io_output_payload_state_elements_10 = io_inputs_2_payload_state_elements_10;
        _zz_io_output_payload_state_elements_11 = io_inputs_2_payload_state_elements_11;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 2'b00) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 2'b01) && io_output_ready);
  assign io_inputs_2_ready = ((io_select == 2'b10) && io_output_ready);
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_round_index = _zz_io_output_payload_round_index;
  assign io_output_payload_state_size = _zz_io_output_payload_state_size;
  assign io_output_payload_state_id = _zz_io_output_payload_state_id;
  assign io_output_payload_state_elements_0 = _zz_io_output_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = _zz_io_output_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = _zz_io_output_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = _zz_io_output_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = _zz_io_output_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = _zz_io_output_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = _zz_io_output_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = _zz_io_output_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = _zz_io_output_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = _zz_io_output_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = _zz_io_output_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = _zz_io_output_payload_state_elements_11;

endmodule

module StreamFifoLowLatency_1 (
  input               io_push_valid,
  output              io_push_ready,
  input      [1:0]    io_push_payload,
  output reg          io_pop_valid,
  input               io_pop_ready,
  output reg [1:0]    io_pop_payload,
  input               io_flush,
  output reg [3:0]    io_occupancy,
  input               clk,
  input               reset
);
  wire       [1:0]    _zz_ram_port0;
  wire       [3:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [3:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  wire       [1:0]    _zz_ram_port;
  wire       [3:0]    _zz_io_occupancy;
  reg                 _zz_1;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [3:0]    pushPtr_valueNext;
  reg        [3:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [3:0]    popPtr_valueNext;
  reg        [3:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                empty;
  wire                full;
  wire                pushing;
  wire                popping;
  wire                when_Stream_l995;
  wire                when_Stream_l1008;
  wire       [3:0]    ptrDif;
  (* ram_style = "distributed" *) reg [1:0] ram [0:8];

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {3'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {3'd0, _zz_popPtr_valueNext_1};
  assign _zz_io_occupancy = (4'b1001 + ptrDif);
  assign _zz_ram_port = io_push_payload;
  assign _zz_ram_port0 = ram[popPtr_value];
  always @(posedge clk) begin
    if(_zz_1) begin
      ram[pushPtr_value] <= _zz_ram_port;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(io_flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 4'b1000);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    if(pushPtr_willOverflow) begin
      pushPtr_valueNext = 4'b0000;
    end else begin
      pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    end
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 4'b0000;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(io_flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 4'b1000);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    if(popPtr_willOverflow) begin
      popPtr_valueNext = 4'b0000;
    end else begin
      popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    end
    if(popPtr_willClear) begin
      popPtr_valueNext = 4'b0000;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign pushing = (io_push_valid && io_push_ready);
  assign popping = (io_pop_valid && io_pop_ready);
  assign io_push_ready = (! full);
  assign when_Stream_l995 = (! empty);
  always @(*) begin
    if(when_Stream_l995) begin
      io_pop_valid = 1'b1;
    end else begin
      io_pop_valid = io_push_valid;
    end
  end

  always @(*) begin
    if(when_Stream_l995) begin
      io_pop_payload = _zz_ram_port0;
    end else begin
      io_pop_payload = io_push_payload;
    end
  end

  assign when_Stream_l1008 = (pushing != popping);
  assign ptrDif = (pushPtr_value - popPtr_value);
  always @(*) begin
    if(ptrMatch) begin
      io_occupancy = (risingOccupancy ? 4'b1001 : 4'b0000);
    end else begin
      io_occupancy = ((popPtr_value < pushPtr_value) ? ptrDif : _zz_io_occupancy);
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      pushPtr_value <= 4'b0000;
      popPtr_value <= 4'b0000;
      risingOccupancy <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      if(when_Stream_l1008) begin
        risingOccupancy <= pushing;
      end
      if(io_flush) begin
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

//StreamDemux replaced by StreamDemux

//StreamFork_10 replaced by StreamFork_10

module MDSMatrixMultiplier_2 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_8 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_9 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_10 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_11 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier_1 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix_4 mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_5 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_6 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_7 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module MDSMatrixMultiplier (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_elements_0,
  output     [254:0]  io_output_payload_state_elements_1,
  output     [254:0]  io_output_payload_state_elements_2,
  output     [254:0]  io_output_payload_state_elements_3,
  output     [254:0]  io_output_payload_state_elements_4,
  output     [254:0]  io_output_payload_state_elements_5,
  output     [254:0]  io_output_payload_state_elements_6,
  output     [254:0]  io_output_payload_state_elements_7,
  output     [254:0]  io_output_payload_state_elements_8,
  output     [254:0]  io_output_payload_state_elements_9,
  output     [254:0]  io_output_payload_state_elements_10,
  output     [254:0]  io_output_payload_state_elements_11,
  input               reset,
  input               clk
);
  wire       [1:0]    mdsMatrix_t3_io_address_port;
  wire       [2:0]    mdsMatrix_t5_io_address_port;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t3_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t5_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t9_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_0;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_1;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_2;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_3;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_4;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_5;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_6;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_7;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_8;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_9;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_10;
  wire       [254:0]  mdsMatrix_t12_io_data_ports_11;
  wire                io_input_translated_fork_io_input_ready;
  wire                io_input_translated_fork_io_outputs_0_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_0_payload;
  wire                io_input_translated_fork_io_outputs_1_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_1_payload;
  wire                io_input_translated_fork_io_outputs_2_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_2_payload;
  wire                io_input_translated_fork_io_outputs_3_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_3_payload;
  wire                io_input_translated_fork_io_outputs_4_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_4_payload;
  wire                io_input_translated_fork_io_outputs_5_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_5_payload;
  wire                io_input_translated_fork_io_outputs_6_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_6_payload;
  wire                io_input_translated_fork_io_outputs_7_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_7_payload;
  wire                io_input_translated_fork_io_outputs_8_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_8_payload;
  wire                io_input_translated_fork_io_outputs_9_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_9_payload;
  wire                io_input_translated_fork_io_outputs_10_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_10_payload;
  wire                io_input_translated_fork_io_outputs_11_valid;
  wire       [254:0]  io_input_translated_fork_io_outputs_11_payload;
  wire                modMultipliers_0_op_ready_o;
  wire                modMultipliers_0_res_valid_o;
  wire       [254:0]  modMultipliers_0_res_o;
  wire                modMultipliers_1_op_ready_o;
  wire                modMultipliers_1_res_valid_o;
  wire       [254:0]  modMultipliers_1_res_o;
  wire                modMultipliers_2_op_ready_o;
  wire                modMultipliers_2_res_valid_o;
  wire       [254:0]  modMultipliers_2_res_o;
  wire                modMultipliers_3_op_ready_o;
  wire                modMultipliers_3_res_valid_o;
  wire       [254:0]  modMultipliers_3_res_o;
  wire                modMultipliers_4_op_ready_o;
  wire                modMultipliers_4_res_valid_o;
  wire       [254:0]  modMultipliers_4_res_o;
  wire                modMultipliers_5_op_ready_o;
  wire                modMultipliers_5_res_valid_o;
  wire       [254:0]  modMultipliers_5_res_o;
  wire                modMultipliers_6_op_ready_o;
  wire                modMultipliers_6_res_valid_o;
  wire       [254:0]  modMultipliers_6_res_o;
  wire                modMultipliers_7_op_ready_o;
  wire                modMultipliers_7_res_valid_o;
  wire       [254:0]  modMultipliers_7_res_o;
  wire                modMultipliers_8_op_ready_o;
  wire                modMultipliers_8_res_valid_o;
  wire       [254:0]  modMultipliers_8_res_o;
  wire                modMultipliers_9_op_ready_o;
  wire                modMultipliers_9_res_valid_o;
  wire       [254:0]  modMultipliers_9_res_o;
  wire                modMultipliers_10_op_ready_o;
  wire                modMultipliers_10_res_valid_o;
  wire       [254:0]  modMultipliers_10_res_o;
  wire                modMultipliers_11_op_ready_o;
  wire                modMultipliers_11_res_valid_o;
  wire       [254:0]  modMultipliers_11_res_o;
  wire       [254:0]  _zz__zz_mulOp2s_0_4;
  wire       [254:0]  _zz__zz_mulOp2s_0_4_1;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  _zz__zz_mulResJoined_translated_payload_state_elements_0_1;
  reg        [254:0]  mulOp2s_0;
  reg        [254:0]  mulOp2s_1;
  reg        [254:0]  mulOp2s_2;
  reg        [254:0]  mulOp2s_3;
  reg        [254:0]  mulOp2s_4;
  reg        [254:0]  mulOp2s_5;
  reg        [254:0]  mulOp2s_6;
  reg        [254:0]  mulOp2s_7;
  reg        [254:0]  mulOp2s_8;
  reg        [254:0]  mulOp2s_9;
  reg        [254:0]  mulOp2s_10;
  reg        [254:0]  mulOp2s_11;
  wire       [3059:0] _zz_mulOp2s_0;
  wire                when_MDSMatrixMultiplier_l51;
  wire       [3059:0] _zz_mulOp2s_0_1;
  wire       [3059:0] _zz_mulOp2s_0_2;
  wire       [3059:0] _zz_mulOp2s_0_3;
  wire       [3059:0] _zz_mulOp2s_0_4;
  wire       [3059:0] _zz_mulOp2s_0_5;
  wire                io_input_translated_valid;
  wire                io_input_translated_ready;
  wire       [254:0]  io_input_translated_payload;
  reg        [6:0]    mulContext_round_index;
  reg        [3:0]    mulContext_state_size;
  reg        [6:0]    mulContext_state_id;
  wire                io_input_fire;
  wire                mulResJoined_valid;
  wire                mulResJoined_ready;
  wire                mulResJoined_fire;
  wire       [3059:0] _zz_mulResJoined_translated_payload_state_elements_0;
  wire                mulResJoined_translated_valid;
  reg                 mulResJoined_translated_ready;
  wire       [6:0]    mulResJoined_translated_payload_round_index;
  wire       [3:0]    mulResJoined_translated_payload_state_size;
  wire       [6:0]    mulResJoined_translated_payload_state_id;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_payload_state_elements_11;
  wire                mulResJoined_translated_m2sPipe_valid;
  wire                mulResJoined_translated_m2sPipe_ready;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_round_index;
  wire       [3:0]    mulResJoined_translated_m2sPipe_payload_state_size;
  wire       [6:0]    mulResJoined_translated_m2sPipe_payload_state_id;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_0;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_1;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_2;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_3;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_4;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_5;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_6;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_7;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_8;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_9;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_10;
  wire       [254:0]  mulResJoined_translated_m2sPipe_payload_state_elements_11;
  reg                 mulResJoined_translated_rValid;
  reg        [6:0]    mulResJoined_translated_rData_round_index;
  reg        [3:0]    mulResJoined_translated_rData_state_size;
  reg        [6:0]    mulResJoined_translated_rData_state_id;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_0;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_1;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_2;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_3;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_4;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_5;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_6;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_7;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_8;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_9;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_10;
  reg        [254:0]  mulResJoined_translated_rData_state_elements_11;
  wire                when_Stream_l342;

  assign _zz__zz_mulOp2s_0_4 = mdsMatrix_t12_io_data_ports_1;
  assign _zz__zz_mulOp2s_0_4_1 = mdsMatrix_t12_io_data_ports_0;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0 = modMultipliers_1_res_o;
  assign _zz__zz_mulResJoined_translated_payload_state_elements_0_1 = modMultipliers_0_res_o;
  MDSMatrix mdsMatrix_t3 (
    .io_data_ports_0    (mdsMatrix_t3_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t3_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t3_io_data_ports_2  ), //o
    .io_address_port    (mdsMatrix_t3_io_address_port  )  //i
  );
  MDSMatrix_1 mdsMatrix_t5 (
    .io_data_ports_0    (mdsMatrix_t5_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t5_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t5_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t5_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t5_io_data_ports_4  ), //o
    .io_address_port    (mdsMatrix_t5_io_address_port  )  //i
  );
  MDSMatrix_2 mdsMatrix_t9 (
    .io_data_ports_0    (mdsMatrix_t9_io_data_ports_0  ), //o
    .io_data_ports_1    (mdsMatrix_t9_io_data_ports_1  ), //o
    .io_data_ports_2    (mdsMatrix_t9_io_data_ports_2  ), //o
    .io_data_ports_3    (mdsMatrix_t9_io_data_ports_3  ), //o
    .io_data_ports_4    (mdsMatrix_t9_io_data_ports_4  ), //o
    .io_data_ports_5    (mdsMatrix_t9_io_data_ports_5  ), //o
    .io_data_ports_6    (mdsMatrix_t9_io_data_ports_6  ), //o
    .io_data_ports_7    (mdsMatrix_t9_io_data_ports_7  ), //o
    .io_data_ports_8    (mdsMatrix_t9_io_data_ports_8  ), //o
    .io_address_port    (io_input_payload_state_index  )  //i
  );
  MDSMatrix_3 mdsMatrix_t12 (
    .io_data_ports_0     (mdsMatrix_t12_io_data_ports_0   ), //o
    .io_data_ports_1     (mdsMatrix_t12_io_data_ports_1   ), //o
    .io_data_ports_2     (mdsMatrix_t12_io_data_ports_2   ), //o
    .io_data_ports_3     (mdsMatrix_t12_io_data_ports_3   ), //o
    .io_data_ports_4     (mdsMatrix_t12_io_data_ports_4   ), //o
    .io_data_ports_5     (mdsMatrix_t12_io_data_ports_5   ), //o
    .io_data_ports_6     (mdsMatrix_t12_io_data_ports_6   ), //o
    .io_data_ports_7     (mdsMatrix_t12_io_data_ports_7   ), //o
    .io_data_ports_8     (mdsMatrix_t12_io_data_ports_8   ), //o
    .io_data_ports_9     (mdsMatrix_t12_io_data_ports_9   ), //o
    .io_data_ports_10    (mdsMatrix_t12_io_data_ports_10  ), //o
    .io_data_ports_11    (mdsMatrix_t12_io_data_ports_11  ), //o
    .io_address_port     (io_input_payload_state_index    )  //i
  );
  StreamFork io_input_translated_fork (
    .io_input_valid           (io_input_translated_valid                       ), //i
    .io_input_ready           (io_input_translated_fork_io_input_ready         ), //o
    .io_input_payload         (io_input_translated_payload                     ), //i
    .io_outputs_0_valid       (io_input_translated_fork_io_outputs_0_valid     ), //o
    .io_outputs_0_ready       (modMultipliers_0_op_ready_o                     ), //i
    .io_outputs_0_payload     (io_input_translated_fork_io_outputs_0_payload   ), //o
    .io_outputs_1_valid       (io_input_translated_fork_io_outputs_1_valid     ), //o
    .io_outputs_1_ready       (modMultipliers_1_op_ready_o                     ), //i
    .io_outputs_1_payload     (io_input_translated_fork_io_outputs_1_payload   ), //o
    .io_outputs_2_valid       (io_input_translated_fork_io_outputs_2_valid     ), //o
    .io_outputs_2_ready       (modMultipliers_2_op_ready_o                     ), //i
    .io_outputs_2_payload     (io_input_translated_fork_io_outputs_2_payload   ), //o
    .io_outputs_3_valid       (io_input_translated_fork_io_outputs_3_valid     ), //o
    .io_outputs_3_ready       (modMultipliers_3_op_ready_o                     ), //i
    .io_outputs_3_payload     (io_input_translated_fork_io_outputs_3_payload   ), //o
    .io_outputs_4_valid       (io_input_translated_fork_io_outputs_4_valid     ), //o
    .io_outputs_4_ready       (modMultipliers_4_op_ready_o                     ), //i
    .io_outputs_4_payload     (io_input_translated_fork_io_outputs_4_payload   ), //o
    .io_outputs_5_valid       (io_input_translated_fork_io_outputs_5_valid     ), //o
    .io_outputs_5_ready       (modMultipliers_5_op_ready_o                     ), //i
    .io_outputs_5_payload     (io_input_translated_fork_io_outputs_5_payload   ), //o
    .io_outputs_6_valid       (io_input_translated_fork_io_outputs_6_valid     ), //o
    .io_outputs_6_ready       (modMultipliers_6_op_ready_o                     ), //i
    .io_outputs_6_payload     (io_input_translated_fork_io_outputs_6_payload   ), //o
    .io_outputs_7_valid       (io_input_translated_fork_io_outputs_7_valid     ), //o
    .io_outputs_7_ready       (modMultipliers_7_op_ready_o                     ), //i
    .io_outputs_7_payload     (io_input_translated_fork_io_outputs_7_payload   ), //o
    .io_outputs_8_valid       (io_input_translated_fork_io_outputs_8_valid     ), //o
    .io_outputs_8_ready       (modMultipliers_8_op_ready_o                     ), //i
    .io_outputs_8_payload     (io_input_translated_fork_io_outputs_8_payload   ), //o
    .io_outputs_9_valid       (io_input_translated_fork_io_outputs_9_valid     ), //o
    .io_outputs_9_ready       (modMultipliers_9_op_ready_o                     ), //i
    .io_outputs_9_payload     (io_input_translated_fork_io_outputs_9_payload   ), //o
    .io_outputs_10_valid      (io_input_translated_fork_io_outputs_10_valid    ), //o
    .io_outputs_10_ready      (modMultipliers_10_op_ready_o                    ), //i
    .io_outputs_10_payload    (io_input_translated_fork_io_outputs_10_payload  ), //o
    .io_outputs_11_valid      (io_input_translated_fork_io_outputs_11_valid    ), //o
    .io_outputs_11_ready      (modMultipliers_11_op_ready_o                    ), //i
    .io_outputs_11_payload    (io_input_translated_fork_io_outputs_11_payload  )  //o
  );
  ModMultiplier modMultipliers_0 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_0_valid    ), //i
    .op_ready_o     (modMultipliers_0_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_0_payload  ), //i
    .op2_i          (mulOp2s_0                                      ), //i
    .res_valid_o    (modMultipliers_0_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_0_res_o                         )  //o
  );
  ModMultiplier modMultipliers_1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_1_valid    ), //i
    .op_ready_o     (modMultipliers_1_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_1_payload  ), //i
    .op2_i          (mulOp2s_1                                      ), //i
    .res_valid_o    (modMultipliers_1_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_1_res_o                         )  //o
  );
  ModMultiplier modMultipliers_2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_2_valid    ), //i
    .op_ready_o     (modMultipliers_2_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_2_payload  ), //i
    .op2_i          (mulOp2s_2                                      ), //i
    .res_valid_o    (modMultipliers_2_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_2_res_o                         )  //o
  );
  ModMultiplier modMultipliers_3 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_3_valid    ), //i
    .op_ready_o     (modMultipliers_3_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_3_payload  ), //i
    .op2_i          (mulOp2s_3                                      ), //i
    .res_valid_o    (modMultipliers_3_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_3_res_o                         )  //o
  );
  ModMultiplier modMultipliers_4 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_4_valid    ), //i
    .op_ready_o     (modMultipliers_4_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_4_payload  ), //i
    .op2_i          (mulOp2s_4                                      ), //i
    .res_valid_o    (modMultipliers_4_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_4_res_o                         )  //o
  );
  ModMultiplier modMultipliers_5 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_5_valid    ), //i
    .op_ready_o     (modMultipliers_5_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_5_payload  ), //i
    .op2_i          (mulOp2s_5                                      ), //i
    .res_valid_o    (modMultipliers_5_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_5_res_o                         )  //o
  );
  ModMultiplier modMultipliers_6 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_6_valid    ), //i
    .op_ready_o     (modMultipliers_6_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_6_payload  ), //i
    .op2_i          (mulOp2s_6                                      ), //i
    .res_valid_o    (modMultipliers_6_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_6_res_o                         )  //o
  );
  ModMultiplier modMultipliers_7 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_7_valid    ), //i
    .op_ready_o     (modMultipliers_7_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_7_payload  ), //i
    .op2_i          (mulOp2s_7                                      ), //i
    .res_valid_o    (modMultipliers_7_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_7_res_o                         )  //o
  );
  ModMultiplier modMultipliers_8 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_8_valid    ), //i
    .op_ready_o     (modMultipliers_8_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_8_payload  ), //i
    .op2_i          (mulOp2s_8                                      ), //i
    .res_valid_o    (modMultipliers_8_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_8_res_o                         )  //o
  );
  ModMultiplier modMultipliers_9 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_9_valid    ), //i
    .op_ready_o     (modMultipliers_9_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_9_payload  ), //i
    .op2_i          (mulOp2s_9                                      ), //i
    .res_valid_o    (modMultipliers_9_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                              ), //i
    .res_o          (modMultipliers_9_res_o                         )  //o
  );
  ModMultiplier modMultipliers_10 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_10_valid    ), //i
    .op_ready_o     (modMultipliers_10_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_10_payload  ), //i
    .op2_i          (mulOp2s_10                                      ), //i
    .res_valid_o    (modMultipliers_10_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_10_res_o                         )  //o
  );
  ModMultiplier modMultipliers_11 (
    .clk            (clk                                             ), //i
    .rst            (reset                                           ), //i
    .op_valid_i     (io_input_translated_fork_io_outputs_11_valid    ), //i
    .op_ready_o     (modMultipliers_11_op_ready_o                    ), //o
    .op1_i          (io_input_translated_fork_io_outputs_11_payload  ), //i
    .op2_i          (mulOp2s_11                                      ), //i
    .res_valid_o    (modMultipliers_11_res_valid_o                   ), //o
    .res_ready_i    (mulResJoined_fire                               ), //i
    .res_o          (modMultipliers_11_res_o                         )  //o
  );
  assign mdsMatrix_t3_io_address_port = io_input_payload_state_index[1:0];
  assign mdsMatrix_t5_io_address_port = io_input_payload_state_index[2:0];
  assign _zz_mulOp2s_0 = {2295'h0,{mdsMatrix_t3_io_data_ports_2,{mdsMatrix_t3_io_data_ports_1,mdsMatrix_t3_io_data_ports_0}}};
  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_0 = _zz_mulOp2s_0[254 : 0];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_0 = _zz_mulOp2s_0_1[254 : 0];
        end else begin
          mulOp2s_0 = _zz_mulOp2s_0_2[254 : 0];
        end
      end
      4'b1001 : begin
        mulOp2s_0 = _zz_mulOp2s_0_3[254 : 0];
      end
      4'b1100 : begin
        mulOp2s_0 = _zz_mulOp2s_0_4[254 : 0];
      end
      default : begin
        mulOp2s_0 = _zz_mulOp2s_0_5[254 : 0];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_1 = _zz_mulOp2s_0[509 : 255];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_1 = _zz_mulOp2s_0_1[509 : 255];
        end else begin
          mulOp2s_1 = _zz_mulOp2s_0_2[509 : 255];
        end
      end
      4'b1001 : begin
        mulOp2s_1 = _zz_mulOp2s_0_3[509 : 255];
      end
      4'b1100 : begin
        mulOp2s_1 = _zz_mulOp2s_0_4[509 : 255];
      end
      default : begin
        mulOp2s_1 = _zz_mulOp2s_0_5[509 : 255];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_2 = _zz_mulOp2s_0[764 : 510];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_2 = _zz_mulOp2s_0_1[764 : 510];
        end else begin
          mulOp2s_2 = _zz_mulOp2s_0_2[764 : 510];
        end
      end
      4'b1001 : begin
        mulOp2s_2 = _zz_mulOp2s_0_3[764 : 510];
      end
      4'b1100 : begin
        mulOp2s_2 = _zz_mulOp2s_0_4[764 : 510];
      end
      default : begin
        mulOp2s_2 = _zz_mulOp2s_0_5[764 : 510];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_3 = _zz_mulOp2s_0[1019 : 765];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_3 = _zz_mulOp2s_0_1[1019 : 765];
        end else begin
          mulOp2s_3 = _zz_mulOp2s_0_2[1019 : 765];
        end
      end
      4'b1001 : begin
        mulOp2s_3 = _zz_mulOp2s_0_3[1019 : 765];
      end
      4'b1100 : begin
        mulOp2s_3 = _zz_mulOp2s_0_4[1019 : 765];
      end
      default : begin
        mulOp2s_3 = _zz_mulOp2s_0_5[1019 : 765];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_4 = _zz_mulOp2s_0[1274 : 1020];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_4 = _zz_mulOp2s_0_1[1274 : 1020];
        end else begin
          mulOp2s_4 = _zz_mulOp2s_0_2[1274 : 1020];
        end
      end
      4'b1001 : begin
        mulOp2s_4 = _zz_mulOp2s_0_3[1274 : 1020];
      end
      4'b1100 : begin
        mulOp2s_4 = _zz_mulOp2s_0_4[1274 : 1020];
      end
      default : begin
        mulOp2s_4 = _zz_mulOp2s_0_5[1274 : 1020];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_5 = _zz_mulOp2s_0[1529 : 1275];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_5 = _zz_mulOp2s_0_1[1529 : 1275];
        end else begin
          mulOp2s_5 = _zz_mulOp2s_0_2[1529 : 1275];
        end
      end
      4'b1001 : begin
        mulOp2s_5 = _zz_mulOp2s_0_3[1529 : 1275];
      end
      4'b1100 : begin
        mulOp2s_5 = _zz_mulOp2s_0_4[1529 : 1275];
      end
      default : begin
        mulOp2s_5 = _zz_mulOp2s_0_5[1529 : 1275];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_6 = _zz_mulOp2s_0[1784 : 1530];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_6 = _zz_mulOp2s_0_1[1784 : 1530];
        end else begin
          mulOp2s_6 = _zz_mulOp2s_0_2[1784 : 1530];
        end
      end
      4'b1001 : begin
        mulOp2s_6 = _zz_mulOp2s_0_3[1784 : 1530];
      end
      4'b1100 : begin
        mulOp2s_6 = _zz_mulOp2s_0_4[1784 : 1530];
      end
      default : begin
        mulOp2s_6 = _zz_mulOp2s_0_5[1784 : 1530];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_7 = _zz_mulOp2s_0[2039 : 1785];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_7 = _zz_mulOp2s_0_1[2039 : 1785];
        end else begin
          mulOp2s_7 = _zz_mulOp2s_0_2[2039 : 1785];
        end
      end
      4'b1001 : begin
        mulOp2s_7 = _zz_mulOp2s_0_3[2039 : 1785];
      end
      4'b1100 : begin
        mulOp2s_7 = _zz_mulOp2s_0_4[2039 : 1785];
      end
      default : begin
        mulOp2s_7 = _zz_mulOp2s_0_5[2039 : 1785];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_8 = _zz_mulOp2s_0[2294 : 2040];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_8 = _zz_mulOp2s_0_1[2294 : 2040];
        end else begin
          mulOp2s_8 = _zz_mulOp2s_0_2[2294 : 2040];
        end
      end
      4'b1001 : begin
        mulOp2s_8 = _zz_mulOp2s_0_3[2294 : 2040];
      end
      4'b1100 : begin
        mulOp2s_8 = _zz_mulOp2s_0_4[2294 : 2040];
      end
      default : begin
        mulOp2s_8 = _zz_mulOp2s_0_5[2294 : 2040];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_9 = _zz_mulOp2s_0[2549 : 2295];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_9 = _zz_mulOp2s_0_1[2549 : 2295];
        end else begin
          mulOp2s_9 = _zz_mulOp2s_0_2[2549 : 2295];
        end
      end
      4'b1001 : begin
        mulOp2s_9 = _zz_mulOp2s_0_3[2549 : 2295];
      end
      4'b1100 : begin
        mulOp2s_9 = _zz_mulOp2s_0_4[2549 : 2295];
      end
      default : begin
        mulOp2s_9 = _zz_mulOp2s_0_5[2549 : 2295];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_10 = _zz_mulOp2s_0[2804 : 2550];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_10 = _zz_mulOp2s_0_1[2804 : 2550];
        end else begin
          mulOp2s_10 = _zz_mulOp2s_0_2[2804 : 2550];
        end
      end
      4'b1001 : begin
        mulOp2s_10 = _zz_mulOp2s_0_3[2804 : 2550];
      end
      4'b1100 : begin
        mulOp2s_10 = _zz_mulOp2s_0_4[2804 : 2550];
      end
      default : begin
        mulOp2s_10 = _zz_mulOp2s_0_5[2804 : 2550];
      end
    endcase
  end

  always @(*) begin
    case(io_input_payload_state_size)
      4'b0011 : begin
        mulOp2s_11 = _zz_mulOp2s_0[3059 : 2805];
      end
      4'b0101 : begin
        if(when_MDSMatrixMultiplier_l51) begin
          mulOp2s_11 = _zz_mulOp2s_0_1[3059 : 2805];
        end else begin
          mulOp2s_11 = _zz_mulOp2s_0_2[3059 : 2805];
        end
      end
      4'b1001 : begin
        mulOp2s_11 = _zz_mulOp2s_0_3[3059 : 2805];
      end
      4'b1100 : begin
        mulOp2s_11 = _zz_mulOp2s_0_4[3059 : 2805];
      end
      default : begin
        mulOp2s_11 = _zz_mulOp2s_0_5[3059 : 2805];
      end
    endcase
  end

  assign when_MDSMatrixMultiplier_l51 = (io_input_payload_state_index == 4'b0101);
  assign _zz_mulOp2s_0_1 = 3060'h0;
  assign _zz_mulOp2s_0_2 = {1785'h0,{mdsMatrix_t5_io_data_ports_4,{mdsMatrix_t5_io_data_ports_3,{mdsMatrix_t5_io_data_ports_2,{mdsMatrix_t5_io_data_ports_1,mdsMatrix_t5_io_data_ports_0}}}}};
  assign _zz_mulOp2s_0_3 = {765'h0,{mdsMatrix_t9_io_data_ports_8,{mdsMatrix_t9_io_data_ports_7,{mdsMatrix_t9_io_data_ports_6,{mdsMatrix_t9_io_data_ports_5,{mdsMatrix_t9_io_data_ports_4,{mdsMatrix_t9_io_data_ports_3,{mdsMatrix_t9_io_data_ports_2,{mdsMatrix_t9_io_data_ports_1,mdsMatrix_t9_io_data_ports_0}}}}}}}}};
  assign _zz_mulOp2s_0_4 = {mdsMatrix_t12_io_data_ports_11,{mdsMatrix_t12_io_data_ports_10,{mdsMatrix_t12_io_data_ports_9,{mdsMatrix_t12_io_data_ports_8,{mdsMatrix_t12_io_data_ports_7,{mdsMatrix_t12_io_data_ports_6,{mdsMatrix_t12_io_data_ports_5,{mdsMatrix_t12_io_data_ports_4,{mdsMatrix_t12_io_data_ports_3,{mdsMatrix_t12_io_data_ports_2,{_zz__zz_mulOp2s_0_4,_zz__zz_mulOp2s_0_4_1}}}}}}}}}}};
  assign _zz_mulOp2s_0_5 = 3060'h0;
  assign io_input_translated_valid = io_input_valid;
  assign io_input_ready = io_input_translated_ready;
  assign io_input_translated_payload = io_input_payload_state_element;
  assign io_input_translated_ready = io_input_translated_fork_io_input_ready;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign mulResJoined_fire = (mulResJoined_valid && mulResJoined_ready);
  assign mulResJoined_valid = (((((((((((modMultipliers_0_res_valid_o && modMultipliers_1_res_valid_o) && modMultipliers_2_res_valid_o) && modMultipliers_3_res_valid_o) && modMultipliers_4_res_valid_o) && modMultipliers_5_res_valid_o) && modMultipliers_6_res_valid_o) && modMultipliers_7_res_valid_o) && modMultipliers_8_res_valid_o) && modMultipliers_9_res_valid_o) && modMultipliers_10_res_valid_o) && modMultipliers_11_res_valid_o);
  assign _zz_mulResJoined_translated_payload_state_elements_0 = {modMultipliers_11_res_o,{modMultipliers_10_res_o,{modMultipliers_9_res_o,{modMultipliers_8_res_o,{modMultipliers_7_res_o,{modMultipliers_6_res_o,{modMultipliers_5_res_o,{modMultipliers_4_res_o,{modMultipliers_3_res_o,{modMultipliers_2_res_o,{_zz__zz_mulResJoined_translated_payload_state_elements_0,_zz__zz_mulResJoined_translated_payload_state_elements_0_1}}}}}}}}}}};
  assign mulResJoined_translated_valid = mulResJoined_valid;
  assign mulResJoined_ready = mulResJoined_translated_ready;
  assign mulResJoined_translated_payload_round_index = mulContext_round_index;
  assign mulResJoined_translated_payload_state_size = mulContext_state_size;
  assign mulResJoined_translated_payload_state_id = mulContext_state_id;
  assign mulResJoined_translated_payload_state_elements_0 = _zz_mulResJoined_translated_payload_state_elements_0[254 : 0];
  assign mulResJoined_translated_payload_state_elements_1 = _zz_mulResJoined_translated_payload_state_elements_0[509 : 255];
  assign mulResJoined_translated_payload_state_elements_2 = _zz_mulResJoined_translated_payload_state_elements_0[764 : 510];
  assign mulResJoined_translated_payload_state_elements_3 = _zz_mulResJoined_translated_payload_state_elements_0[1019 : 765];
  assign mulResJoined_translated_payload_state_elements_4 = _zz_mulResJoined_translated_payload_state_elements_0[1274 : 1020];
  assign mulResJoined_translated_payload_state_elements_5 = _zz_mulResJoined_translated_payload_state_elements_0[1529 : 1275];
  assign mulResJoined_translated_payload_state_elements_6 = _zz_mulResJoined_translated_payload_state_elements_0[1784 : 1530];
  assign mulResJoined_translated_payload_state_elements_7 = _zz_mulResJoined_translated_payload_state_elements_0[2039 : 1785];
  assign mulResJoined_translated_payload_state_elements_8 = _zz_mulResJoined_translated_payload_state_elements_0[2294 : 2040];
  assign mulResJoined_translated_payload_state_elements_9 = _zz_mulResJoined_translated_payload_state_elements_0[2549 : 2295];
  assign mulResJoined_translated_payload_state_elements_10 = _zz_mulResJoined_translated_payload_state_elements_0[2804 : 2550];
  assign mulResJoined_translated_payload_state_elements_11 = _zz_mulResJoined_translated_payload_state_elements_0[3059 : 2805];
  always @(*) begin
    mulResJoined_translated_ready = mulResJoined_translated_m2sPipe_ready;
    if(when_Stream_l342) begin
      mulResJoined_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mulResJoined_translated_m2sPipe_valid);
  assign mulResJoined_translated_m2sPipe_valid = mulResJoined_translated_rValid;
  assign mulResJoined_translated_m2sPipe_payload_round_index = mulResJoined_translated_rData_round_index;
  assign mulResJoined_translated_m2sPipe_payload_state_size = mulResJoined_translated_rData_state_size;
  assign mulResJoined_translated_m2sPipe_payload_state_id = mulResJoined_translated_rData_state_id;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_0 = mulResJoined_translated_rData_state_elements_0;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_1 = mulResJoined_translated_rData_state_elements_1;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_2 = mulResJoined_translated_rData_state_elements_2;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_3 = mulResJoined_translated_rData_state_elements_3;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_4 = mulResJoined_translated_rData_state_elements_4;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_5 = mulResJoined_translated_rData_state_elements_5;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_6 = mulResJoined_translated_rData_state_elements_6;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_7 = mulResJoined_translated_rData_state_elements_7;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_8 = mulResJoined_translated_rData_state_elements_8;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_9 = mulResJoined_translated_rData_state_elements_9;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_10 = mulResJoined_translated_rData_state_elements_10;
  assign mulResJoined_translated_m2sPipe_payload_state_elements_11 = mulResJoined_translated_rData_state_elements_11;
  assign io_output_valid = mulResJoined_translated_m2sPipe_valid;
  assign mulResJoined_translated_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mulResJoined_translated_m2sPipe_payload_round_index;
  assign io_output_payload_state_size = mulResJoined_translated_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mulResJoined_translated_m2sPipe_payload_state_id;
  assign io_output_payload_state_elements_0 = mulResJoined_translated_m2sPipe_payload_state_elements_0;
  assign io_output_payload_state_elements_1 = mulResJoined_translated_m2sPipe_payload_state_elements_1;
  assign io_output_payload_state_elements_2 = mulResJoined_translated_m2sPipe_payload_state_elements_2;
  assign io_output_payload_state_elements_3 = mulResJoined_translated_m2sPipe_payload_state_elements_3;
  assign io_output_payload_state_elements_4 = mulResJoined_translated_m2sPipe_payload_state_elements_4;
  assign io_output_payload_state_elements_5 = mulResJoined_translated_m2sPipe_payload_state_elements_5;
  assign io_output_payload_state_elements_6 = mulResJoined_translated_m2sPipe_payload_state_elements_6;
  assign io_output_payload_state_elements_7 = mulResJoined_translated_m2sPipe_payload_state_elements_7;
  assign io_output_payload_state_elements_8 = mulResJoined_translated_m2sPipe_payload_state_elements_8;
  assign io_output_payload_state_elements_9 = mulResJoined_translated_m2sPipe_payload_state_elements_9;
  assign io_output_payload_state_elements_10 = mulResJoined_translated_m2sPipe_payload_state_elements_10;
  assign io_output_payload_state_elements_11 = mulResJoined_translated_m2sPipe_payload_state_elements_11;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mulContext_state_size <= 4'b0000;
      mulContext_state_id <= 7'h0;
      mulContext_round_index <= 7'h0;
      mulResJoined_translated_rValid <= 1'b0;
    end else begin
      if(io_input_fire) begin
        mulContext_round_index <= io_input_payload_round_index;
        mulContext_state_size <= io_input_payload_state_size;
        mulContext_state_id <= io_input_payload_state_id;
      end
      if(mulResJoined_translated_ready) begin
        mulResJoined_translated_rValid <= mulResJoined_translated_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mulResJoined_translated_ready) begin
      mulResJoined_translated_rData_round_index <= mulResJoined_translated_payload_round_index;
      mulResJoined_translated_rData_state_size <= mulResJoined_translated_payload_state_size;
      mulResJoined_translated_rData_state_id <= mulResJoined_translated_payload_state_id;
      mulResJoined_translated_rData_state_elements_0 <= mulResJoined_translated_payload_state_elements_0;
      mulResJoined_translated_rData_state_elements_1 <= mulResJoined_translated_payload_state_elements_1;
      mulResJoined_translated_rData_state_elements_2 <= mulResJoined_translated_payload_state_elements_2;
      mulResJoined_translated_rData_state_elements_3 <= mulResJoined_translated_payload_state_elements_3;
      mulResJoined_translated_rData_state_elements_4 <= mulResJoined_translated_payload_state_elements_4;
      mulResJoined_translated_rData_state_elements_5 <= mulResJoined_translated_payload_state_elements_5;
      mulResJoined_translated_rData_state_elements_6 <= mulResJoined_translated_payload_state_elements_6;
      mulResJoined_translated_rData_state_elements_7 <= mulResJoined_translated_payload_state_elements_7;
      mulResJoined_translated_rData_state_elements_8 <= mulResJoined_translated_payload_state_elements_8;
      mulResJoined_translated_rData_state_elements_9 <= mulResJoined_translated_payload_state_elements_9;
      mulResJoined_translated_rData_state_elements_10 <= mulResJoined_translated_payload_state_elements_10;
      mulResJoined_translated_rData_state_elements_11 <= mulResJoined_translated_payload_state_elements_11;
    end
  end


endmodule

module StreamMux (
  input      [1:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [6:0]    io_inputs_0_payload_round_index,
  input      [3:0]    io_inputs_0_payload_state_index,
  input      [3:0]    io_inputs_0_payload_state_size,
  input      [6:0]    io_inputs_0_payload_state_id,
  input      [254:0]  io_inputs_0_payload_state_element,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [6:0]    io_inputs_1_payload_round_index,
  input      [3:0]    io_inputs_1_payload_state_index,
  input      [3:0]    io_inputs_1_payload_state_size,
  input      [6:0]    io_inputs_1_payload_state_id,
  input      [254:0]  io_inputs_1_payload_state_element,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [6:0]    io_inputs_2_payload_round_index,
  input      [3:0]    io_inputs_2_payload_state_index,
  input      [3:0]    io_inputs_2_payload_state_size,
  input      [6:0]    io_inputs_2_payload_state_id,
  input      [254:0]  io_inputs_2_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_element
);
  reg                 _zz_io_output_valid;
  reg        [6:0]    _zz_io_output_payload_round_index;
  reg        [3:0]    _zz_io_output_payload_state_index;
  reg        [3:0]    _zz_io_output_payload_state_size;
  reg        [6:0]    _zz_io_output_payload_state_id;
  reg        [254:0]  _zz_io_output_payload_state_element;

  always @(*) begin
    case(io_select)
      2'b00 : begin
        _zz_io_output_valid = io_inputs_0_valid;
        _zz_io_output_payload_round_index = io_inputs_0_payload_round_index;
        _zz_io_output_payload_state_index = io_inputs_0_payload_state_index;
        _zz_io_output_payload_state_size = io_inputs_0_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_0_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_0_payload_state_element;
      end
      2'b01 : begin
        _zz_io_output_valid = io_inputs_1_valid;
        _zz_io_output_payload_round_index = io_inputs_1_payload_round_index;
        _zz_io_output_payload_state_index = io_inputs_1_payload_state_index;
        _zz_io_output_payload_state_size = io_inputs_1_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_1_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_1_payload_state_element;
      end
      default : begin
        _zz_io_output_valid = io_inputs_2_valid;
        _zz_io_output_payload_round_index = io_inputs_2_payload_round_index;
        _zz_io_output_payload_state_index = io_inputs_2_payload_state_index;
        _zz_io_output_payload_state_size = io_inputs_2_payload_state_size;
        _zz_io_output_payload_state_id = io_inputs_2_payload_state_id;
        _zz_io_output_payload_state_element = io_inputs_2_payload_state_element;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 2'b00) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 2'b01) && io_output_ready);
  assign io_inputs_2_ready = ((io_select == 2'b10) && io_output_ready);
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_round_index = _zz_io_output_payload_round_index;
  assign io_output_payload_state_index = _zz_io_output_payload_state_index;
  assign io_output_payload_state_size = _zz_io_output_payload_state_size;
  assign io_output_payload_state_id = _zz_io_output_payload_state_id;
  assign io_output_payload_state_element = _zz_io_output_payload_state_element;

endmodule

module StreamFifoLowLatency (
  input               io_push_valid,
  output              io_push_ready,
  input      [1:0]    io_push_payload,
  output reg          io_pop_valid,
  input               io_pop_ready,
  output reg [1:0]    io_pop_payload,
  input               io_flush,
  output reg [4:0]    io_occupancy,
  input               clk,
  input               reset
);
  wire       [1:0]    _zz_ram_port0;
  wire       [4:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [4:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  wire       [1:0]    _zz_ram_port;
  wire       [4:0]    _zz_io_occupancy;
  reg                 _zz_1;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [4:0]    pushPtr_valueNext;
  reg        [4:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [4:0]    popPtr_valueNext;
  reg        [4:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                empty;
  wire                full;
  wire                pushing;
  wire                popping;
  wire                when_Stream_l995;
  wire                when_Stream_l1008;
  wire       [4:0]    ptrDif;
  (* ram_style = "distributed" *) reg [1:0] ram [0:19];

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {4'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {4'd0, _zz_popPtr_valueNext_1};
  assign _zz_io_occupancy = (5'h14 + ptrDif);
  assign _zz_ram_port = io_push_payload;
  assign _zz_ram_port0 = ram[popPtr_value];
  always @(posedge clk) begin
    if(_zz_1) begin
      ram[pushPtr_value] <= _zz_ram_port;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(io_flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 5'h13);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    if(pushPtr_willOverflow) begin
      pushPtr_valueNext = 5'h0;
    end else begin
      pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    end
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 5'h0;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(io_flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 5'h13);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    if(popPtr_willOverflow) begin
      popPtr_valueNext = 5'h0;
    end else begin
      popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    end
    if(popPtr_willClear) begin
      popPtr_valueNext = 5'h0;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign pushing = (io_push_valid && io_push_ready);
  assign popping = (io_pop_valid && io_pop_ready);
  assign io_push_ready = (! full);
  assign when_Stream_l995 = (! empty);
  always @(*) begin
    if(when_Stream_l995) begin
      io_pop_valid = 1'b1;
    end else begin
      io_pop_valid = io_push_valid;
    end
  end

  always @(*) begin
    if(when_Stream_l995) begin
      io_pop_payload = _zz_ram_port0;
    end else begin
      io_pop_payload = io_push_payload;
    end
  end

  assign when_Stream_l1008 = (pushing != popping);
  assign ptrDif = (pushPtr_value - popPtr_value);
  always @(*) begin
    if(ptrMatch) begin
      io_occupancy = (risingOccupancy ? 5'h14 : 5'h0);
    end else begin
      io_occupancy = ((popPtr_value < pushPtr_value) ? ptrDif : _zz_io_occupancy);
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      pushPtr_value <= 5'h0;
      popPtr_value <= 5'h0;
      risingOccupancy <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      if(when_Stream_l1008) begin
        risingOccupancy <= pushing;
      end
      if(io_flush) begin
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamDemux (
  input      [1:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_round_index,
  output     [3:0]    io_outputs_0_payload_state_index,
  output     [3:0]    io_outputs_0_payload_state_size,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [254:0]  io_outputs_0_payload_state_element,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_round_index,
  output     [3:0]    io_outputs_1_payload_state_index,
  output     [3:0]    io_outputs_1_payload_state_size,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [254:0]  io_outputs_1_payload_state_element,
  output reg          io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [6:0]    io_outputs_2_payload_round_index,
  output     [3:0]    io_outputs_2_payload_state_index,
  output     [3:0]    io_outputs_2_payload_state_size,
  output     [6:0]    io_outputs_2_payload_state_id,
  output     [254:0]  io_outputs_2_payload_state_element
);
  wire                when_Stream_l745;
  wire                when_Stream_l745_1;
  wire                when_Stream_l745_2;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l745) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l745_1) begin
      io_input_ready = io_outputs_1_ready;
    end
    if(!when_Stream_l745_2) begin
      io_input_ready = io_outputs_2_ready;
    end
  end

  assign io_outputs_0_payload_round_index = io_input_payload_round_index;
  assign io_outputs_0_payload_state_index = io_input_payload_state_index;
  assign io_outputs_0_payload_state_size = io_input_payload_state_size;
  assign io_outputs_0_payload_state_id = io_input_payload_state_id;
  assign io_outputs_0_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745 = (2'b00 != io_select);
  always @(*) begin
    if(when_Stream_l745) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_round_index = io_input_payload_round_index;
  assign io_outputs_1_payload_state_index = io_input_payload_state_index;
  assign io_outputs_1_payload_state_size = io_input_payload_state_size;
  assign io_outputs_1_payload_state_id = io_input_payload_state_id;
  assign io_outputs_1_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_1 = (2'b01 != io_select);
  always @(*) begin
    if(when_Stream_l745_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end

  assign io_outputs_2_payload_round_index = io_input_payload_round_index;
  assign io_outputs_2_payload_state_index = io_input_payload_state_index;
  assign io_outputs_2_payload_state_size = io_input_payload_state_size;
  assign io_outputs_2_payload_state_id = io_input_payload_state_id;
  assign io_outputs_2_payload_state_element = io_input_payload_state_element;
  assign when_Stream_l745_2 = (2'b10 != io_select);
  always @(*) begin
    if(when_Stream_l745_2) begin
      io_outputs_2_valid = 1'b0;
    end else begin
      io_outputs_2_valid = io_input_valid;
    end
  end


endmodule

module StreamFork_10 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_round_index,
  output     [3:0]    io_outputs_0_payload_state_index,
  output     [3:0]    io_outputs_0_payload_state_size,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [254:0]  io_outputs_0_payload_state_element,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_round_index,
  output     [3:0]    io_outputs_1_payload_state_index,
  output     [3:0]    io_outputs_1_payload_state_size,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [254:0]  io_outputs_1_payload_state_element
);

  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_round_index = io_input_payload_round_index;
  assign io_outputs_0_payload_state_index = io_input_payload_state_index;
  assign io_outputs_0_payload_state_size = io_input_payload_state_size;
  assign io_outputs_0_payload_state_id = io_input_payload_state_id;
  assign io_outputs_0_payload_state_element = io_input_payload_state_element;
  assign io_outputs_1_payload_round_index = io_input_payload_round_index;
  assign io_outputs_1_payload_state_index = io_input_payload_state_index;
  assign io_outputs_1_payload_state_size = io_input_payload_state_size;
  assign io_outputs_1_payload_state_id = io_input_payload_state_id;
  assign io_outputs_1_payload_state_element = io_input_payload_state_element;

endmodule

//SBox5 replaced by SBox5

//SBox5 replaced by SBox5

module SBox5 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [254:0]  io_input_payload_state_element,
  output              io_output_valid,
  input               io_output_ready,
  output     [6:0]    io_output_payload_round_index,
  output     [3:0]    io_output_payload_state_index,
  output     [3:0]    io_output_payload_state_size,
  output     [6:0]    io_output_payload_state_id,
  output     [254:0]  io_output_payload_state_element,
  input               reset,
  input               clk
);
  wire                mul_stage0_multiplier0_op_ready_o;
  wire                mul_stage0_multiplier0_res_valid_o;
  wire       [254:0]  mul_stage0_multiplier0_res_o;
  wire                mul_stage1_multiplier1_op_ready_o;
  wire                mul_stage1_multiplier1_res_valid_o;
  wire       [254:0]  mul_stage1_multiplier1_res_o;
  wire                mul_stage2_multiplier2_op_ready_o;
  wire                mul_stage2_multiplier2_res_valid_o;
  wire       [254:0]  mul_stage2_multiplier2_res_o;
  reg        [6:0]    mul_stage0_mulContext_round_index;
  reg        [3:0]    mul_stage0_mulContext_state_index;
  reg        [3:0]    mul_stage0_mulContext_state_size;
  reg        [6:0]    mul_stage0_mulContext_state_id;
  reg        [254:0]  mul_stage0_mulContext_initial_state;
  wire                mul_stage0_output_valid;
  reg                 mul_stage0_output_ready;
  wire       [6:0]    mul_stage0_output_payload_round_index;
  wire       [3:0]    mul_stage0_output_payload_state_index;
  wire       [3:0]    mul_stage0_output_payload_state_size;
  wire       [6:0]    mul_stage0_output_payload_state_id;
  wire       [254:0]  mul_stage0_output_payload_state_element;
  wire       [254:0]  mul_stage0_output_payload_initial_state;
  wire                mul_stage0_multiplier0_cmd_fire;
  wire                mul_stage0_output_input_valid;
  wire                mul_stage0_output_input_ready;
  wire       [6:0]    mul_stage0_output_input_payload_round_index;
  wire       [3:0]    mul_stage0_output_input_payload_state_index;
  wire       [3:0]    mul_stage0_output_input_payload_state_size;
  wire       [6:0]    mul_stage0_output_input_payload_state_id;
  wire       [254:0]  mul_stage0_output_input_payload_state_element;
  wire       [254:0]  mul_stage0_output_input_payload_initial_state;
  reg                 mul_stage0_output_rValid;
  reg        [6:0]    mul_stage0_output_rData_round_index;
  reg        [3:0]    mul_stage0_output_rData_state_index;
  reg        [3:0]    mul_stage0_output_rData_state_size;
  reg        [6:0]    mul_stage0_output_rData_state_id;
  reg        [254:0]  mul_stage0_output_rData_state_element;
  reg        [254:0]  mul_stage0_output_rData_initial_state;
  wire                when_Stream_l342;
  reg        [6:0]    mul_stage1_mulContext_round_index;
  reg        [3:0]    mul_stage1_mulContext_state_index;
  reg        [3:0]    mul_stage1_mulContext_state_size;
  reg        [6:0]    mul_stage1_mulContext_state_id;
  reg        [254:0]  mul_stage1_mulContext_initial_state;
  wire                mul_stage1_output_valid;
  reg                 mul_stage1_output_ready;
  wire       [6:0]    mul_stage1_output_payload_round_index;
  wire       [3:0]    mul_stage1_output_payload_state_index;
  wire       [3:0]    mul_stage1_output_payload_state_size;
  wire       [6:0]    mul_stage1_output_payload_state_id;
  wire       [254:0]  mul_stage1_output_payload_state_element;
  wire       [254:0]  mul_stage1_output_payload_initial_state;
  wire                mul_stage1_multiplier1_cmd_fire;
  wire                mul_stage1_output_input_valid;
  wire                mul_stage1_output_input_ready;
  wire       [6:0]    mul_stage1_output_input_payload_round_index;
  wire       [3:0]    mul_stage1_output_input_payload_state_index;
  wire       [3:0]    mul_stage1_output_input_payload_state_size;
  wire       [6:0]    mul_stage1_output_input_payload_state_id;
  wire       [254:0]  mul_stage1_output_input_payload_state_element;
  wire       [254:0]  mul_stage1_output_input_payload_initial_state;
  reg                 mul_stage1_output_rValid;
  reg        [6:0]    mul_stage1_output_rData_round_index;
  reg        [3:0]    mul_stage1_output_rData_state_index;
  reg        [3:0]    mul_stage1_output_rData_state_size;
  reg        [6:0]    mul_stage1_output_rData_state_id;
  reg        [254:0]  mul_stage1_output_rData_state_element;
  reg        [254:0]  mul_stage1_output_rData_initial_state;
  wire                when_Stream_l342_1;
  reg        [6:0]    mul_stage2_mulContext_round_index;
  reg        [3:0]    mul_stage2_mulContext_state_index;
  reg        [3:0]    mul_stage2_mulContext_state_size;
  reg        [6:0]    mul_stage2_mulContext_state_id;
  reg        [254:0]  mul_stage2_mulContext_initial_state;
  wire                mul_stage2_output_valid;
  reg                 mul_stage2_output_ready;
  wire       [6:0]    mul_stage2_output_payload_round_index;
  wire       [3:0]    mul_stage2_output_payload_state_index;
  wire       [3:0]    mul_stage2_output_payload_state_size;
  wire       [6:0]    mul_stage2_output_payload_state_id;
  wire       [254:0]  mul_stage2_output_payload_state_element;
  wire                mul_stage2_multiplier2_cmd_fire;
  reg                 mul_stage2_is_partial_round;
  wire                mul_stage2_is_pass_sbox5;
  wire                mul_stage2_output_m2sPipe_valid;
  wire                mul_stage2_output_m2sPipe_ready;
  wire       [6:0]    mul_stage2_output_m2sPipe_payload_round_index;
  wire       [3:0]    mul_stage2_output_m2sPipe_payload_state_index;
  wire       [3:0]    mul_stage2_output_m2sPipe_payload_state_size;
  wire       [6:0]    mul_stage2_output_m2sPipe_payload_state_id;
  wire       [254:0]  mul_stage2_output_m2sPipe_payload_state_element;
  reg                 mul_stage2_output_rValid;
  reg        [6:0]    mul_stage2_output_rData_round_index;
  reg        [3:0]    mul_stage2_output_rData_state_index;
  reg        [3:0]    mul_stage2_output_rData_state_size;
  reg        [6:0]    mul_stage2_output_rData_state_id;
  reg        [254:0]  mul_stage2_output_rData_state_element;
  wire                when_Stream_l342_2;

  ModMultiplier mul_stage0_multiplier0 (
    .clk            (clk                                 ), //i
    .rst            (reset                               ), //i
    .op_valid_i     (io_input_valid                      ), //i
    .op_ready_o     (mul_stage0_multiplier0_op_ready_o   ), //o
    .op1_i          (io_input_payload_state_element      ), //i
    .op2_i          (io_input_payload_state_element      ), //i
    .res_valid_o    (mul_stage0_multiplier0_res_valid_o  ), //o
    .res_ready_i    (mul_stage0_output_ready             ), //i
    .res_o          (mul_stage0_multiplier0_res_o        )  //o
  );
  ModMultiplier mul_stage1_multiplier1 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (mul_stage0_output_input_valid                  ), //i
    .op_ready_o     (mul_stage1_multiplier1_op_ready_o              ), //o
    .op1_i          (mul_stage0_output_input_payload_state_element  ), //i
    .op2_i          (mul_stage0_output_input_payload_state_element  ), //i
    .res_valid_o    (mul_stage1_multiplier1_res_valid_o             ), //o
    .res_ready_i    (mul_stage1_output_ready                        ), //i
    .res_o          (mul_stage1_multiplier1_res_o                   )  //o
  );
  ModMultiplier mul_stage2_multiplier2 (
    .clk            (clk                                            ), //i
    .rst            (reset                                          ), //i
    .op_valid_i     (mul_stage1_output_input_valid                  ), //i
    .op_ready_o     (mul_stage2_multiplier2_op_ready_o              ), //o
    .op1_i          (mul_stage1_output_input_payload_initial_state  ), //i
    .op2_i          (mul_stage1_output_input_payload_state_element  ), //i
    .res_valid_o    (mul_stage2_multiplier2_res_valid_o             ), //o
    .res_ready_i    (mul_stage2_output_ready                        ), //i
    .res_o          (mul_stage2_multiplier2_res_o                   )  //o
  );
  assign io_input_ready = mul_stage0_multiplier0_op_ready_o;
  assign mul_stage0_multiplier0_cmd_fire = (io_input_valid && mul_stage0_multiplier0_op_ready_o);
  assign mul_stage0_output_valid = mul_stage0_multiplier0_res_valid_o;
  assign mul_stage0_output_payload_round_index = mul_stage0_mulContext_round_index;
  assign mul_stage0_output_payload_state_index = mul_stage0_mulContext_state_index;
  assign mul_stage0_output_payload_state_size = mul_stage0_mulContext_state_size;
  assign mul_stage0_output_payload_state_id = mul_stage0_mulContext_state_id;
  assign mul_stage0_output_payload_initial_state = mul_stage0_mulContext_initial_state;
  assign mul_stage0_output_payload_state_element = mul_stage0_multiplier0_res_o;
  always @(*) begin
    mul_stage0_output_ready = mul_stage0_output_input_ready;
    if(when_Stream_l342) begin
      mul_stage0_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! mul_stage0_output_input_valid);
  assign mul_stage0_output_input_valid = mul_stage0_output_rValid;
  assign mul_stage0_output_input_payload_round_index = mul_stage0_output_rData_round_index;
  assign mul_stage0_output_input_payload_state_index = mul_stage0_output_rData_state_index;
  assign mul_stage0_output_input_payload_state_size = mul_stage0_output_rData_state_size;
  assign mul_stage0_output_input_payload_state_id = mul_stage0_output_rData_state_id;
  assign mul_stage0_output_input_payload_state_element = mul_stage0_output_rData_state_element;
  assign mul_stage0_output_input_payload_initial_state = mul_stage0_output_rData_initial_state;
  assign mul_stage0_output_input_ready = mul_stage1_multiplier1_op_ready_o;
  assign mul_stage1_multiplier1_cmd_fire = (mul_stage0_output_input_valid && mul_stage1_multiplier1_op_ready_o);
  assign mul_stage1_output_valid = mul_stage1_multiplier1_res_valid_o;
  assign mul_stage1_output_payload_round_index = mul_stage1_mulContext_round_index;
  assign mul_stage1_output_payload_state_index = mul_stage1_mulContext_state_index;
  assign mul_stage1_output_payload_state_size = mul_stage1_mulContext_state_size;
  assign mul_stage1_output_payload_state_id = mul_stage1_mulContext_state_id;
  assign mul_stage1_output_payload_initial_state = mul_stage1_mulContext_initial_state;
  assign mul_stage1_output_payload_state_element = mul_stage1_multiplier1_res_o;
  always @(*) begin
    mul_stage1_output_ready = mul_stage1_output_input_ready;
    if(when_Stream_l342_1) begin
      mul_stage1_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! mul_stage1_output_input_valid);
  assign mul_stage1_output_input_valid = mul_stage1_output_rValid;
  assign mul_stage1_output_input_payload_round_index = mul_stage1_output_rData_round_index;
  assign mul_stage1_output_input_payload_state_index = mul_stage1_output_rData_state_index;
  assign mul_stage1_output_input_payload_state_size = mul_stage1_output_rData_state_size;
  assign mul_stage1_output_input_payload_state_id = mul_stage1_output_rData_state_id;
  assign mul_stage1_output_input_payload_state_element = mul_stage1_output_rData_state_element;
  assign mul_stage1_output_input_payload_initial_state = mul_stage1_output_rData_initial_state;
  assign mul_stage1_output_input_ready = mul_stage2_multiplier2_op_ready_o;
  assign mul_stage2_multiplier2_cmd_fire = (mul_stage1_output_input_valid && mul_stage2_multiplier2_op_ready_o);
  assign mul_stage2_output_valid = mul_stage2_multiplier2_res_valid_o;
  assign mul_stage2_output_payload_round_index = mul_stage2_mulContext_round_index;
  assign mul_stage2_output_payload_state_index = mul_stage2_mulContext_state_index;
  assign mul_stage2_output_payload_state_size = mul_stage2_mulContext_state_size;
  assign mul_stage2_output_payload_state_id = mul_stage2_mulContext_state_id;
  always @(*) begin
    case(mul_stage2_mulContext_state_size)
      4'b0011 : begin
        mul_stage2_is_partial_round = ((7'h04 <= mul_stage2_mulContext_round_index) && (mul_stage2_mulContext_round_index < 7'h3b));
      end
      4'b0101 : begin
        mul_stage2_is_partial_round = ((7'h04 <= mul_stage2_mulContext_round_index) && (mul_stage2_mulContext_round_index < 7'h3c));
      end
      4'b1001 : begin
        mul_stage2_is_partial_round = ((7'h04 <= mul_stage2_mulContext_round_index) && (mul_stage2_mulContext_round_index < 7'h3d));
      end
      4'b1100 : begin
        mul_stage2_is_partial_round = ((7'h04 <= mul_stage2_mulContext_round_index) && (mul_stage2_mulContext_round_index < 7'h3d));
      end
      default : begin
        mul_stage2_is_partial_round = 1'b0;
      end
    endcase
  end

  assign mul_stage2_is_pass_sbox5 = (mul_stage2_is_partial_round && (mul_stage2_mulContext_state_index != 4'b0000));
  assign mul_stage2_output_payload_state_element = (mul_stage2_is_pass_sbox5 ? mul_stage2_mulContext_initial_state : mul_stage2_multiplier2_res_o);
  always @(*) begin
    mul_stage2_output_ready = mul_stage2_output_m2sPipe_ready;
    if(when_Stream_l342_2) begin
      mul_stage2_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342_2 = (! mul_stage2_output_m2sPipe_valid);
  assign mul_stage2_output_m2sPipe_valid = mul_stage2_output_rValid;
  assign mul_stage2_output_m2sPipe_payload_round_index = mul_stage2_output_rData_round_index;
  assign mul_stage2_output_m2sPipe_payload_state_index = mul_stage2_output_rData_state_index;
  assign mul_stage2_output_m2sPipe_payload_state_size = mul_stage2_output_rData_state_size;
  assign mul_stage2_output_m2sPipe_payload_state_id = mul_stage2_output_rData_state_id;
  assign mul_stage2_output_m2sPipe_payload_state_element = mul_stage2_output_rData_state_element;
  assign io_output_valid = mul_stage2_output_m2sPipe_valid;
  assign mul_stage2_output_m2sPipe_ready = io_output_ready;
  assign io_output_payload_round_index = mul_stage2_output_m2sPipe_payload_round_index;
  assign io_output_payload_state_index = mul_stage2_output_m2sPipe_payload_state_index;
  assign io_output_payload_state_size = mul_stage2_output_m2sPipe_payload_state_size;
  assign io_output_payload_state_id = mul_stage2_output_m2sPipe_payload_state_id;
  assign io_output_payload_state_element = mul_stage2_output_m2sPipe_payload_state_element;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mul_stage0_mulContext_state_index <= 4'b0000;
      mul_stage0_mulContext_round_index <= 7'h0;
      mul_stage0_mulContext_state_size <= 4'b0000;
      mul_stage0_mulContext_initial_state <= 255'h0;
      mul_stage0_output_rValid <= 1'b0;
      mul_stage1_mulContext_state_index <= 4'b0000;
      mul_stage1_mulContext_round_index <= 7'h0;
      mul_stage1_mulContext_state_size <= 4'b0000;
      mul_stage1_mulContext_initial_state <= 255'h0;
      mul_stage1_output_rValid <= 1'b0;
      mul_stage2_mulContext_state_index <= 4'b0000;
      mul_stage2_mulContext_round_index <= 7'h0;
      mul_stage2_mulContext_state_size <= 4'b0000;
      mul_stage2_mulContext_initial_state <= 255'h0;
      mul_stage2_output_rValid <= 1'b0;
    end else begin
      if(mul_stage0_multiplier0_cmd_fire) begin
        mul_stage0_mulContext_round_index <= io_input_payload_round_index;
        mul_stage0_mulContext_state_index <= io_input_payload_state_index;
        mul_stage0_mulContext_state_size <= io_input_payload_state_size;
        mul_stage0_mulContext_initial_state <= io_input_payload_state_element;
      end
      if(mul_stage0_output_ready) begin
        mul_stage0_output_rValid <= mul_stage0_output_valid;
      end
      if(mul_stage1_multiplier1_cmd_fire) begin
        mul_stage1_mulContext_round_index <= mul_stage0_output_input_payload_round_index;
        mul_stage1_mulContext_state_index <= mul_stage0_output_input_payload_state_index;
        mul_stage1_mulContext_state_size <= mul_stage0_output_input_payload_state_size;
        mul_stage1_mulContext_initial_state <= mul_stage0_output_input_payload_initial_state;
      end
      if(mul_stage1_output_ready) begin
        mul_stage1_output_rValid <= mul_stage1_output_valid;
      end
      if(mul_stage2_multiplier2_cmd_fire) begin
        mul_stage2_mulContext_round_index <= mul_stage1_output_input_payload_round_index;
        mul_stage2_mulContext_state_index <= mul_stage1_output_input_payload_state_index;
        mul_stage2_mulContext_state_size <= mul_stage1_output_input_payload_state_size;
        mul_stage2_mulContext_initial_state <= mul_stage1_output_input_payload_initial_state;
      end
      if(mul_stage2_output_ready) begin
        mul_stage2_output_rValid <= mul_stage2_output_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(mul_stage0_multiplier0_cmd_fire) begin
      mul_stage0_mulContext_state_id <= io_input_payload_state_id;
    end
    if(mul_stage0_output_ready) begin
      mul_stage0_output_rData_round_index <= mul_stage0_output_payload_round_index;
      mul_stage0_output_rData_state_index <= mul_stage0_output_payload_state_index;
      mul_stage0_output_rData_state_size <= mul_stage0_output_payload_state_size;
      mul_stage0_output_rData_state_id <= mul_stage0_output_payload_state_id;
      mul_stage0_output_rData_state_element <= mul_stage0_output_payload_state_element;
      mul_stage0_output_rData_initial_state <= mul_stage0_output_payload_initial_state;
    end
    if(mul_stage1_multiplier1_cmd_fire) begin
      mul_stage1_mulContext_state_id <= mul_stage0_output_input_payload_state_id;
    end
    if(mul_stage1_output_ready) begin
      mul_stage1_output_rData_round_index <= mul_stage1_output_payload_round_index;
      mul_stage1_output_rData_state_index <= mul_stage1_output_payload_state_index;
      mul_stage1_output_rData_state_size <= mul_stage1_output_payload_state_size;
      mul_stage1_output_rData_state_id <= mul_stage1_output_payload_state_id;
      mul_stage1_output_rData_state_element <= mul_stage1_output_payload_state_element;
      mul_stage1_output_rData_initial_state <= mul_stage1_output_payload_initial_state;
    end
    if(mul_stage2_multiplier2_cmd_fire) begin
      mul_stage2_mulContext_state_id <= mul_stage1_output_input_payload_state_id;
    end
    if(mul_stage2_output_ready) begin
      mul_stage2_output_rData_round_index <= mul_stage2_output_payload_round_index;
      mul_stage2_output_rData_state_index <= mul_stage2_output_payload_state_index;
      mul_stage2_output_rData_state_size <= mul_stage2_output_payload_state_size;
      mul_stage2_output_rData_state_id <= mul_stage2_output_payload_state_id;
      mul_stage2_output_rData_state_element <= mul_stage2_output_payload_state_element;
    end
  end


endmodule

module RoundConstants_3 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  wire       [254:0]  _zz_constants_roms_9_port0;
  wire       [254:0]  _zz_constants_roms_10_port0;
  wire       [254:0]  _zz_constants_roms_11_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_9 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_10 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_11 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_9.bin",constants_roms_9);
  end
  assign _zz_constants_roms_9_port0 = constants_roms_9[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_10.bin",constants_roms_10);
  end
  assign _zz_constants_roms_10_port0 = constants_roms_10[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t12_constants_roms_11.bin",constants_roms_11);
  end
  assign _zz_constants_roms_11_port0 = constants_roms_11[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      4'b1000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
      4'b1001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_9_port0;
      end
      4'b1010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_10_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_11_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_2 (
  output     [254:0]  io_read_ports_0_data,
  input      [3:0]    io_read_ports_0_t_index,
  input      [6:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  wire       [254:0]  _zz_constants_roms_5_port0;
  wire       [254:0]  _zz_constants_roms_6_port0;
  wire       [254:0]  _zz_constants_roms_7_port0;
  wire       [254:0]  _zz_constants_roms_8_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_5 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_6 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_7 [0:64];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_8 [0:64];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_5.bin",constants_roms_5);
  end
  assign _zz_constants_roms_5_port0 = constants_roms_5[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_6.bin",constants_roms_6);
  end
  assign _zz_constants_roms_6_port0 = constants_roms_6[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_7.bin",constants_roms_7);
  end
  assign _zz_constants_roms_7_port0 = constants_roms_7[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t9_constants_roms_8.bin",constants_roms_8);
  end
  assign _zz_constants_roms_8_port0 = constants_roms_8[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      4'b0000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      4'b0001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      4'b0010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      4'b0011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      4'b0100 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
      4'b0101 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_5_port0;
      end
      4'b0110 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_6_port0;
      end
      4'b0111 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_7_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_8_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants_1 (
  output     [254:0]  io_read_ports_0_data,
  input      [2:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  wire       [254:0]  _zz_constants_roms_3_port0;
  wire       [254:0]  _zz_constants_roms_4_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_3 [0:63];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_4 [0:63];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t5_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t5_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t5_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t5_constants_roms_3.bin",constants_roms_3);
  end
  assign _zz_constants_roms_3_port0 = constants_roms_3[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t5_constants_roms_4.bin",constants_roms_4);
  end
  assign _zz_constants_roms_4_port0 = constants_roms_4[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      3'b000 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      3'b001 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      3'b010 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
      3'b011 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_3_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_4_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module RoundConstants (
  output     [254:0]  io_read_ports_0_data,
  input      [1:0]    io_read_ports_0_t_index,
  input      [5:0]    io_read_ports_0_round_index
);
  wire       [254:0]  _zz_constants_roms_0_port0;
  wire       [254:0]  _zz_constants_roms_1_port0;
  wire       [254:0]  _zz_constants_roms_2_port0;
  reg        [254:0]  _zz_io_read_ports_0_data;
  (* ram_style = "distributed" *) reg [254:0] constants_roms_0 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_1 [0:62];
  (* ram_style = "distributed" *) reg [254:0] constants_roms_2 [0:62];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t3_constants_roms_0.bin",constants_roms_0);
  end
  assign _zz_constants_roms_0_port0 = constants_roms_0[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t3_constants_roms_1.bin",constants_roms_1);
  end
  assign _zz_constants_roms_1_port0 = constants_roms_1[io_read_ports_0_round_index];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_AddRoundConstantStage_roundConstants_t3_constants_roms_2.bin",constants_roms_2);
  end
  assign _zz_constants_roms_2_port0 = constants_roms_2[io_read_ports_0_round_index];
  always @(*) begin
    case(io_read_ports_0_t_index)
      2'b00 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_0_port0;
      end
      2'b01 : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_1_port0;
      end
      default : begin
        _zz_io_read_ports_0_data = _zz_constants_roms_2_port0;
      end
    endcase
  end

  assign io_read_ports_0_data = _zz_io_read_ports_0_data;

endmodule

module StreamFork_9 (
  input               io_input_valid,
  output              io_input_ready,
  input      [6:0]    io_input_payload_round_index,
  input      [3:0]    io_input_payload_state_size,
  input      [6:0]    io_input_payload_state_id,
  input      [3:0]    io_input_payload_state_indexes_0,
  input      [3:0]    io_input_payload_state_indexes_1,
  input      [3:0]    io_input_payload_state_indexes_2,
  input      [254:0]  io_input_payload_state_elements_0,
  input      [254:0]  io_input_payload_state_elements_1,
  input      [254:0]  io_input_payload_state_elements_2,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [6:0]    io_outputs_0_payload_round_index,
  output     [3:0]    io_outputs_0_payload_state_size,
  output     [6:0]    io_outputs_0_payload_state_id,
  output     [3:0]    io_outputs_0_payload_state_indexes_0,
  output     [3:0]    io_outputs_0_payload_state_indexes_1,
  output     [3:0]    io_outputs_0_payload_state_indexes_2,
  output     [254:0]  io_outputs_0_payload_state_elements_0,
  output     [254:0]  io_outputs_0_payload_state_elements_1,
  output     [254:0]  io_outputs_0_payload_state_elements_2,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [6:0]    io_outputs_1_payload_round_index,
  output     [3:0]    io_outputs_1_payload_state_size,
  output     [6:0]    io_outputs_1_payload_state_id,
  output     [3:0]    io_outputs_1_payload_state_indexes_0,
  output     [3:0]    io_outputs_1_payload_state_indexes_1,
  output     [3:0]    io_outputs_1_payload_state_indexes_2,
  output     [254:0]  io_outputs_1_payload_state_elements_0,
  output     [254:0]  io_outputs_1_payload_state_elements_1,
  output     [254:0]  io_outputs_1_payload_state_elements_2,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [6:0]    io_outputs_2_payload_round_index,
  output     [3:0]    io_outputs_2_payload_state_size,
  output     [6:0]    io_outputs_2_payload_state_id,
  output     [3:0]    io_outputs_2_payload_state_indexes_0,
  output     [3:0]    io_outputs_2_payload_state_indexes_1,
  output     [3:0]    io_outputs_2_payload_state_indexes_2,
  output     [254:0]  io_outputs_2_payload_state_elements_0,
  output     [254:0]  io_outputs_2_payload_state_elements_1,
  output     [254:0]  io_outputs_2_payload_state_elements_2
);

  assign io_input_ready = ((io_outputs_0_ready && io_outputs_1_ready) && io_outputs_2_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_2_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_round_index = io_input_payload_round_index;
  assign io_outputs_0_payload_state_size = io_input_payload_state_size;
  assign io_outputs_0_payload_state_id = io_input_payload_state_id;
  assign io_outputs_0_payload_state_indexes_0 = io_input_payload_state_indexes_0;
  assign io_outputs_0_payload_state_indexes_1 = io_input_payload_state_indexes_1;
  assign io_outputs_0_payload_state_indexes_2 = io_input_payload_state_indexes_2;
  assign io_outputs_0_payload_state_elements_0 = io_input_payload_state_elements_0;
  assign io_outputs_0_payload_state_elements_1 = io_input_payload_state_elements_1;
  assign io_outputs_0_payload_state_elements_2 = io_input_payload_state_elements_2;
  assign io_outputs_1_payload_round_index = io_input_payload_round_index;
  assign io_outputs_1_payload_state_size = io_input_payload_state_size;
  assign io_outputs_1_payload_state_id = io_input_payload_state_id;
  assign io_outputs_1_payload_state_indexes_0 = io_input_payload_state_indexes_0;
  assign io_outputs_1_payload_state_indexes_1 = io_input_payload_state_indexes_1;
  assign io_outputs_1_payload_state_indexes_2 = io_input_payload_state_indexes_2;
  assign io_outputs_1_payload_state_elements_0 = io_input_payload_state_elements_0;
  assign io_outputs_1_payload_state_elements_1 = io_input_payload_state_elements_1;
  assign io_outputs_1_payload_state_elements_2 = io_input_payload_state_elements_2;
  assign io_outputs_2_payload_round_index = io_input_payload_round_index;
  assign io_outputs_2_payload_state_size = io_input_payload_state_size;
  assign io_outputs_2_payload_state_id = io_input_payload_state_id;
  assign io_outputs_2_payload_state_indexes_0 = io_input_payload_state_indexes_0;
  assign io_outputs_2_payload_state_indexes_1 = io_input_payload_state_indexes_1;
  assign io_outputs_2_payload_state_indexes_2 = io_input_payload_state_indexes_2;
  assign io_outputs_2_payload_state_elements_0 = io_input_payload_state_elements_0;
  assign io_outputs_2_payload_state_elements_1 = io_input_payload_state_elements_1;
  assign io_outputs_2_payload_state_elements_2 = io_input_payload_state_elements_2;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_35 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_34 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_33 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_32 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_31 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_30 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_29 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_28 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_27 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_26 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_25 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_24 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_5_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_23 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_22 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_21 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_20 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_19 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_18 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_17 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_16 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_15 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_14 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_13 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_12 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_4_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_11 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_10 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_9 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_8 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_2_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

//StreamFork replaced by StreamFork

module MDSMatrix_7 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_6 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_5 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix_4 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_1_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule

module StreamFork (
  input               io_input_valid,
  output              io_input_ready,
  input      [254:0]  io_input_payload,
  output              io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [254:0]  io_outputs_0_payload,
  output              io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [254:0]  io_outputs_1_payload,
  output              io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [254:0]  io_outputs_2_payload,
  output              io_outputs_3_valid,
  input               io_outputs_3_ready,
  output     [254:0]  io_outputs_3_payload,
  output              io_outputs_4_valid,
  input               io_outputs_4_ready,
  output     [254:0]  io_outputs_4_payload,
  output              io_outputs_5_valid,
  input               io_outputs_5_ready,
  output     [254:0]  io_outputs_5_payload,
  output              io_outputs_6_valid,
  input               io_outputs_6_ready,
  output     [254:0]  io_outputs_6_payload,
  output              io_outputs_7_valid,
  input               io_outputs_7_ready,
  output     [254:0]  io_outputs_7_payload,
  output              io_outputs_8_valid,
  input               io_outputs_8_ready,
  output     [254:0]  io_outputs_8_payload,
  output              io_outputs_9_valid,
  input               io_outputs_9_ready,
  output     [254:0]  io_outputs_9_payload,
  output              io_outputs_10_valid,
  input               io_outputs_10_ready,
  output     [254:0]  io_outputs_10_payload,
  output              io_outputs_11_valid,
  input               io_outputs_11_ready,
  output     [254:0]  io_outputs_11_payload
);

  assign io_input_ready = (((((((((((io_outputs_0_ready && io_outputs_1_ready) && io_outputs_2_ready) && io_outputs_3_ready) && io_outputs_4_ready) && io_outputs_5_ready) && io_outputs_6_ready) && io_outputs_7_ready) && io_outputs_8_ready) && io_outputs_9_ready) && io_outputs_10_ready) && io_outputs_11_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_2_valid = (io_input_valid && io_input_ready);
  assign io_outputs_3_valid = (io_input_valid && io_input_ready);
  assign io_outputs_4_valid = (io_input_valid && io_input_ready);
  assign io_outputs_5_valid = (io_input_valid && io_input_ready);
  assign io_outputs_6_valid = (io_input_valid && io_input_ready);
  assign io_outputs_7_valid = (io_input_valid && io_input_ready);
  assign io_outputs_8_valid = (io_input_valid && io_input_ready);
  assign io_outputs_9_valid = (io_input_valid && io_input_ready);
  assign io_outputs_10_valid = (io_input_valid && io_input_ready);
  assign io_outputs_11_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload = io_input_payload;
  assign io_outputs_1_payload = io_input_payload;
  assign io_outputs_2_payload = io_input_payload;
  assign io_outputs_3_payload = io_input_payload;
  assign io_outputs_4_payload = io_input_payload;
  assign io_outputs_5_payload = io_input_payload;
  assign io_outputs_6_payload = io_input_payload;
  assign io_outputs_7_payload = io_input_payload;
  assign io_outputs_8_payload = io_input_payload;
  assign io_outputs_9_payload = io_input_payload;
  assign io_outputs_10_payload = io_input_payload;
  assign io_outputs_11_payload = io_input_payload;

endmodule

module MDSMatrix_3 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  output     [254:0]  io_data_ports_9,
  output     [254:0]  io_data_ports_10,
  output     [254:0]  io_data_ports_11,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  wire       [254:0]  _zz_mds_roms_9_port0;
  wire       [254:0]  _zz_mds_roms_10_port0;
  wire       [254:0]  _zz_mds_roms_11_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_9 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_10 [0:11];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_11 [0:11];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_9.bin",mds_roms_9);
  end
  assign _zz_mds_roms_9_port0 = mds_roms_9[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_10.bin",mds_roms_10);
  end
  assign _zz_mds_roms_10_port0 = mds_roms_10[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t12_mds_roms_11.bin",mds_roms_11);
  end
  assign _zz_mds_roms_11_port0 = mds_roms_11[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;
  assign io_data_ports_9 = _zz_mds_roms_9_port0;
  assign io_data_ports_10 = _zz_mds_roms_10_port0;
  assign io_data_ports_11 = _zz_mds_roms_11_port0;

endmodule

module MDSMatrix_2 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  output     [254:0]  io_data_ports_5,
  output     [254:0]  io_data_ports_6,
  output     [254:0]  io_data_ports_7,
  output     [254:0]  io_data_ports_8,
  input      [3:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  wire       [254:0]  _zz_mds_roms_5_port0;
  wire       [254:0]  _zz_mds_roms_6_port0;
  wire       [254:0]  _zz_mds_roms_7_port0;
  wire       [254:0]  _zz_mds_roms_8_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_5 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_6 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_7 [0:8];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_8 [0:8];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_5.bin",mds_roms_5);
  end
  assign _zz_mds_roms_5_port0 = mds_roms_5[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_6.bin",mds_roms_6);
  end
  assign _zz_mds_roms_6_port0 = mds_roms_6[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_7.bin",mds_roms_7);
  end
  assign _zz_mds_roms_7_port0 = mds_roms_7[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t9_mds_roms_8.bin",mds_roms_8);
  end
  assign _zz_mds_roms_8_port0 = mds_roms_8[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;
  assign io_data_ports_5 = _zz_mds_roms_5_port0;
  assign io_data_ports_6 = _zz_mds_roms_6_port0;
  assign io_data_ports_7 = _zz_mds_roms_7_port0;
  assign io_data_ports_8 = _zz_mds_roms_8_port0;

endmodule

module MDSMatrix_1 (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  output     [254:0]  io_data_ports_3,
  output     [254:0]  io_data_ports_4,
  input      [2:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  wire       [254:0]  _zz_mds_roms_3_port0;
  wire       [254:0]  _zz_mds_roms_4_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_3 [0:4];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_4 [0:4];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_3.bin",mds_roms_3);
  end
  assign _zz_mds_roms_3_port0 = mds_roms_3[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t5_mds_roms_4.bin",mds_roms_4);
  end
  assign _zz_mds_roms_4_port0 = mds_roms_4[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;
  assign io_data_ports_3 = _zz_mds_roms_3_port0;
  assign io_data_ports_4 = _zz_mds_roms_4_port0;

endmodule

module MDSMatrix (
  output     [254:0]  io_data_ports_0,
  output     [254:0]  io_data_ports_1,
  output     [254:0]  io_data_ports_2,
  input      [1:0]    io_address_port
);
  wire       [254:0]  _zz_mds_roms_0_port0;
  wire       [254:0]  _zz_mds_roms_1_port0;
  wire       [254:0]  _zz_mds_roms_2_port0;
  (* ram_style = "distributed" *) reg [254:0] mds_roms_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_1 [0:2];
  (* ram_style = "distributed" *) reg [254:0] mds_roms_2 [0:2];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_0.bin",mds_roms_0);
  end
  assign _zz_mds_roms_0_port0 = mds_roms_0[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_1.bin",mds_roms_1);
  end
  assign _zz_mds_roms_1_port0 = mds_roms_1[io_address_port];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonThread_3_MDSMixStage_matrixMultiplierInsts_0_mdsMatrix_t3_mds_roms_2.bin",mds_roms_2);
  end
  assign _zz_mds_roms_2_port0 = mds_roms_2[io_address_port];
  assign io_data_ports_0 = _zz_mds_roms_0_port0;
  assign io_data_ports_1 = _zz_mds_roms_1_port0;
  assign io_data_ports_2 = _zz_mds_roms_2_port0;

endmodule
